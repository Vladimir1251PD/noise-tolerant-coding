`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:00:04 05/02/2024 
// Design Name: 
// Module Name:    RAM 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
parameter RAM_WIDTH = 24;
parameter RAM_ADDR_BITS = 12;
module RAM(
	input clk,
	input [RAM_ADDR_BITS-1:0] address,
	output reg [RAM_WIDTH-1:0] output_reg
	
    );

   
   (* RAM_STYLE="{AUTO | BLOCK |  BLOCK_POWER1 | BLOCK_POWER2}" *)
   reg [RAM_WIDTH-1:0] block_ram [(2**RAM_ADDR_BITS)-1:0];

   //  The forllowing code is only necessary if you wish to initialize the RAM 
   //  contents via an external file (use $readmemb for binary data)
   initial
	begin
		output_reg = 0;
      block_ram[0] = 24'b000000000000000000000000 ; 
		block_ram[1] = 24'b000000000000000000000001 ; 
		block_ram[2] = 24'b000000000000000000000010 ; 
		block_ram[3] = 24'b000000000000000000000011 ; 
		block_ram[4] = 24'b000000000000000000000100 ; 
		block_ram[5] = 24'b000000000000000000000101 ; 
		block_ram[6] = 24'b000000000000000000000110 ; 
		block_ram[7] = 24'b000000000000000000000111 ; 
		block_ram[8] = 24'b000000000000000000001000 ; 
		block_ram[9] = 24'b000000000000000000001001 ; 
		block_ram[10] = 24'b000000000000000000001010 ; 
		block_ram[11] = 24'b000000000000000000001011 ; 
		block_ram[12] = 24'b000000000000000000001100 ; 
		block_ram[13] = 24'b000000000000000000001101 ; 
		block_ram[14] = 24'b000000000000000000001110 ; 
		block_ram[15] = 24'b000000000000000000001111 ; 
		block_ram[16] = 24'b000000000000000000010000 ; 
		block_ram[17] = 24'b000000000000000000010001 ; 
		block_ram[18] = 24'b000000000000000000010010 ; 
		block_ram[19] = 24'b000000000000000000010011 ; 
		block_ram[20] = 24'b000000000000000000010100 ; 
		block_ram[21] = 24'b000000000000000000010101 ; 
		block_ram[22] = 24'b000000000000000000010110 ; 
		block_ram[23] = 24'b000000000000000000010111 ; 
		block_ram[24] = 24'b000000000000000000011000 ; 
		block_ram[25] = 24'b000000000000000000011001 ; 
		block_ram[26] = 24'b000000000000000000011010 ; 
		block_ram[27] = 24'b000000000000000000011011 ; 
		block_ram[28] = 24'b000000000000000000011100 ; 
		block_ram[29] = 24'b000000000000000000011101 ; 
		block_ram[30] = 24'b000000000000000000011110 ; 
		block_ram[31] = 24'b010010000000001000000000 ; 
		block_ram[32] = 24'b000000000000000000100000 ; 
		block_ram[33] = 24'b000000000000000000100001 ; 
		block_ram[34] = 24'b000000000000000000100010 ; 
		block_ram[35] = 24'b000000000000000000100011 ; 
		block_ram[36] = 24'b000000000000000000100100 ; 
		block_ram[37] = 24'b000000000000000000100101 ; 
		block_ram[38] = 24'b000000000000000000100110 ; 
		block_ram[39] = 24'b000000000000000000100111 ; 
		block_ram[40] = 24'b000000000000000000101000 ; 
		block_ram[41] = 24'b000000000000000000101001 ; 
		block_ram[42] = 24'b000000000000000000101010 ; 
		block_ram[43] = 24'b000000000000000000101011 ; 
		block_ram[44] = 24'b000000000000000000101100 ; 
		block_ram[45] = 24'b000000000000000000101101 ; 
		block_ram[46] = 24'b000000000000000000101110 ; 
		block_ram[47] = 24'b000000100101000000000000 ; 
		block_ram[48] = 24'b000000000000000000110000 ; 
		block_ram[49] = 24'b000000000000000000110001 ; 
		block_ram[50] = 24'b000000000000000000110010 ; 
		block_ram[51] = 24'b000000000000000000110011 ; 
		block_ram[52] = 24'b000000000000000000110100 ; 
		block_ram[53] = 24'b000000000000000000110101 ; 
		block_ram[54] = 24'b000000000000000000110110 ; 
		block_ram[55] = 24'b000001000000100010000000 ; 
		block_ram[56] = 24'b000000000000000000111000 ; 
		block_ram[57] = 24'b000000000000000000111001 ; 
		block_ram[58] = 24'b000000000000000000111010 ; 
		block_ram[59] = 24'b000000011000000100000000 ; 
		block_ram[60] = 24'b000000000000000000111100 ; 
		block_ram[61] = 24'b001000000010000001000000 ; 
		block_ram[62] = 24'b100100000000010000000000 ; 
		block_ram[63] = 24'b000000011000000100000100 ; 
		block_ram[64] = 24'b000000000000000001000000 ; 
		block_ram[65] = 24'b000000000000000001000001 ; 
		block_ram[66] = 24'b000000000000000001000010 ; 
		block_ram[67] = 24'b000000000000000001000011 ; 
		block_ram[68] = 24'b000000000000000001000100 ; 
		block_ram[69] = 24'b000000000000000001000101 ; 
		block_ram[70] = 24'b000000000000000001000110 ; 
		block_ram[71] = 24'b000000000000000001000111 ; 
		block_ram[72] = 24'b000000000000000001001000 ; 
		block_ram[73] = 24'b000000000000000001001001 ; 
		block_ram[74] = 24'b000000000000000001001010 ; 
		block_ram[75] = 24'b000000000000000001001011 ; 
		block_ram[76] = 24'b000000000000000001001100 ; 
		block_ram[77] = 24'b000000000000000001001101 ; 
		block_ram[78] = 24'b000000000000000001001110 ; 
		block_ram[79] = 24'b100000010000000010000000 ; 
		block_ram[80] = 24'b000000000000000001010000 ; 
		block_ram[81] = 24'b000000000000000001010001 ; 
		block_ram[82] = 24'b000000000000000001010010 ; 
		block_ram[83] = 24'b000000000000000001010011 ; 
		block_ram[84] = 24'b000000000000000001010100 ; 
		block_ram[85] = 24'b000000000000000001010101 ; 
		block_ram[86] = 24'b000000000000000001010110 ; 
		block_ram[87] = 24'b000100000100000100000000 ; 
		block_ram[88] = 24'b000000000000000001011000 ; 
		block_ram[89] = 24'b000000000000000001011001 ; 
		block_ram[90] = 24'b000000000000000001011010 ; 
		block_ram[91] = 24'b000000100000110000000000 ; 
		block_ram[92] = 24'b000000000000000001011100 ; 
		block_ram[93] = 24'b001000000010000000100000 ; 
		block_ram[94] = 24'b000001001001000000000000 ; 
		block_ram[95] = 24'b000000100000110000000100 ; 
		block_ram[96] = 24'b000000000000000001100000 ; 
		block_ram[97] = 24'b000000000000000001100001 ; 
		block_ram[98] = 24'b000000000000000001100010 ; 
		block_ram[99] = 24'b000000000000000001100011 ; 
		block_ram[100] = 24'b000000000000000001100100 ; 
		block_ram[101] = 24'b000000000000000001100101 ; 
		block_ram[102] = 24'b000000000000000001100110 ; 
		block_ram[103] = 24'b010000001000010000000000 ; 
		block_ram[104] = 24'b000000000000000001101000 ; 
		block_ram[105] = 24'b000000000000000001101001 ; 
		block_ram[106] = 24'b000000000000000001101010 ; 
		block_ram[107] = 24'b000101000000001000000000 ; 
		block_ram[108] = 24'b000000000000000001101100 ; 
		block_ram[109] = 24'b001000000010000000010000 ; 
		block_ram[110] = 24'b000010000000100100000000 ; 
		block_ram[111] = 24'b000000100101000001000000 ; 
		block_ram[112] = 24'b000000000000000001110000 ; 
		block_ram[113] = 24'b000000000000000001110001 ; 
		block_ram[114] = 24'b000000000000000001110010 ; 
		block_ram[115] = 24'b100010000001000000000000 ; 
		block_ram[116] = 24'b000000000000000001110100 ; 
		block_ram[117] = 24'b001000000010000000001000 ; 
		block_ram[118] = 24'b000000110000001000000000 ; 
		block_ram[119] = 24'b000000110000001000000001 ; 
		block_ram[120] = 24'b000000000000000001111000 ; 
		block_ram[121] = 24'b001000000010000000000100 ; 
		block_ram[122] = 24'b010000000100000010000000 ; 
		block_ram[123] = 24'b000000011000000101000000 ; 
		block_ram[124] = 24'b001000000010000000000001 ; 
		block_ram[125] = 24'b001000000010000000000000 ; 
		block_ram[126] = 24'b000000110000001000001000 ; 
		block_ram[127] = 24'b001000000010000000000010 ; 
		block_ram[128] = 24'b000000000000000010000000 ; 
		block_ram[129] = 24'b000000000000000010000001 ; 
		block_ram[130] = 24'b000000000000000010000010 ; 
		block_ram[131] = 24'b000000000000000010000011 ; 
		block_ram[132] = 24'b000000000000000010000100 ; 
		block_ram[133] = 24'b000000000000000010000101 ; 
		block_ram[134] = 24'b000000000000000010000110 ; 
		block_ram[135] = 24'b000000000000000010000111 ; 
		block_ram[136] = 24'b000000000000000010001000 ; 
		block_ram[137] = 24'b000000000000000010001001 ; 
		block_ram[138] = 24'b000000000000000010001010 ; 
		block_ram[139] = 24'b000000000000000010001011 ; 
		block_ram[140] = 24'b000000000000000010001100 ; 
		block_ram[141] = 24'b000000000000000010001101 ; 
		block_ram[142] = 24'b000000000000000010001110 ; 
		block_ram[143] = 24'b100000010000000001000000 ; 
		block_ram[144] = 24'b000000000000000010010000 ; 
		block_ram[145] = 24'b000000000000000010010001 ; 
		block_ram[146] = 24'b000000000000000010010010 ; 
		block_ram[147] = 24'b000000000000000010010011 ; 
		block_ram[148] = 24'b000000000000000010010100 ; 
		block_ram[149] = 24'b000000000000000010010101 ; 
		block_ram[150] = 24'b000000000000000010010110 ; 
		block_ram[151] = 24'b000001000000100000100000 ; 
		block_ram[152] = 24'b000000000000000010011000 ; 
		block_ram[153] = 24'b000000000000000010011001 ; 
		block_ram[154] = 24'b000000000000000010011010 ; 
		block_ram[155] = 24'b001100000001000000000000 ; 
		block_ram[156] = 24'b000000000000000010011100 ; 
		block_ram[157] = 24'b000000001100010000000000 ; 
		block_ram[158] = 24'b000000100010000100000000 ; 
		block_ram[159] = 24'b000000001100010000000010 ; 
		block_ram[160] = 24'b000000000000000010100000 ; 
		block_ram[161] = 24'b000000000000000010100001 ; 
		block_ram[162] = 24'b000000000000000010100010 ; 
		block_ram[163] = 24'b000000000000000010100011 ; 
		block_ram[164] = 24'b000000000000000010100100 ; 
		block_ram[165] = 24'b000000000000000010100101 ; 
		block_ram[166] = 24'b000000000000000010100110 ; 
		block_ram[167] = 24'b000001000000100000010000 ; 
		block_ram[168] = 24'b000000000000000010101000 ; 
		block_ram[169] = 24'b000000000000000010101001 ; 
		block_ram[170] = 24'b000000000000000010101010 ; 
		block_ram[171] = 24'b000010000010010000000000 ; 
		block_ram[172] = 24'b000000000000000010101100 ; 
		block_ram[173] = 24'b010100000000000100000000 ; 
		block_ram[174] = 24'b001000001000001000000000 ; 
		block_ram[175] = 24'b000000100101000010000000 ; 
		block_ram[176] = 24'b000000000000000010110000 ; 
		block_ram[177] = 24'b000000000000000010110001 ; 
		block_ram[178] = 24'b000000000000000010110010 ; 
		block_ram[179] = 24'b000001000000100000000100 ; 
		block_ram[180] = 24'b000000000000000010110100 ; 
		block_ram[181] = 24'b000001000000100000000010 ; 
		block_ram[182] = 24'b000001000000100000000001 ; 
		block_ram[183] = 24'b000001000000100000000000 ; 
		block_ram[184] = 24'b000000000000000010111000 ; 
		block_ram[185] = 24'b100000100000001000000000 ; 
		block_ram[186] = 24'b010000000100000001000000 ; 
		block_ram[187] = 24'b000000011000000110000000 ; 
		block_ram[188] = 24'b000010010001000000000000 ; 
		block_ram[189] = 24'b000000001100010000100000 ; 
		block_ram[190] = 24'b000000100010000100100000 ; 
		block_ram[191] = 24'b000001000000100000001000 ; 
		block_ram[192] = 24'b000000000000000011000000 ; 
		block_ram[193] = 24'b000000000000000011000001 ; 
		block_ram[194] = 24'b000000000000000011000010 ; 
		block_ram[195] = 24'b000000000000000011000011 ; 
		block_ram[196] = 24'b000000000000000011000100 ; 
		block_ram[197] = 24'b000000000000000011000101 ; 
		block_ram[198] = 24'b000000000000000011000110 ; 
		block_ram[199] = 24'b100000010000000000001000 ; 
		block_ram[200] = 24'b000000000000000011001000 ; 
		block_ram[201] = 24'b000000000000000011001001 ; 
		block_ram[202] = 24'b000000000000000011001010 ; 
		block_ram[203] = 24'b100000010000000000000100 ; 
		block_ram[204] = 24'b000000000000000011001100 ; 
		block_ram[205] = 24'b100000010000000000000010 ; 
		block_ram[206] = 24'b100000010000000000000001 ; 
		block_ram[207] = 24'b100000010000000000000000 ; 
		block_ram[208] = 24'b000000000000000011010000 ; 
		block_ram[209] = 24'b000000000000000011010001 ; 
		block_ram[210] = 24'b000000000000000011010010 ; 
		block_ram[211] = 24'b000000001010001000000000 ; 
		block_ram[212] = 24'b000000000000000011010100 ; 
		block_ram[213] = 24'b010000100001000000000000 ; 
		block_ram[214] = 24'b001010000000010000000000 ; 
		block_ram[215] = 24'b000000001010001000000100 ; 
		block_ram[216] = 24'b000000000000000011011000 ; 
		block_ram[217] = 24'b000011000000000100000000 ; 
		block_ram[218] = 24'b010000000100000000100000 ; 
		block_ram[219] = 24'b000000001010001000001000 ; 
		block_ram[220] = 24'b000100000000101000000000 ; 
		block_ram[221] = 24'b000000001100010001000000 ; 
		block_ram[222] = 24'b000000100010000101000000 ; 
		block_ram[223] = 24'b100000010000000000010000 ; 
		block_ram[224] = 24'b000000000000000011100000 ; 
		block_ram[225] = 24'b000000000000000011100001 ; 
		block_ram[226] = 24'b000000000000000011100010 ; 
		block_ram[227] = 24'b001000100000000100000000 ; 
		block_ram[228] = 24'b000000000000000011100100 ; 
		block_ram[229] = 24'b000010000100001000000000 ; 
		block_ram[230] = 24'b000100000011000000000000 ; 
		block_ram[231] = 24'b000001000000100001010000 ; 
		block_ram[232] = 24'b000000000000000011101000 ; 
		block_ram[233] = 24'b000000001001100000000000 ; 
		block_ram[234] = 24'b010000000100000000010000 ; 
		block_ram[235] = 24'b000000001001100000000010 ; 
		block_ram[236] = 24'b000001100000010000000000 ; 
		block_ram[237] = 24'b000000001001100000000100 ; 
		block_ram[238] = 24'b000001100000010000000010 ; 
		block_ram[239] = 24'b100000010000000000100000 ; 
		block_ram[240] = 24'b000000000000000011110000 ; 
		block_ram[241] = 24'b000100010000010000000000 ; 
		block_ram[242] = 24'b010000000100000000001000 ; 
		block_ram[243] = 24'b000000001010001000100000 ; 
		block_ram[244] = 24'b100000001000000100000000 ; 
		block_ram[245] = 24'b000001000000100001000010 ; 
		block_ram[246] = 24'b000000110000001010000000 ; 
		block_ram[247] = 24'b000001000000100001000000 ; 
		block_ram[248] = 24'b010000000100000000000010 ; 
		block_ram[249] = 24'b000000001001100000010000 ; 
		block_ram[250] = 24'b010000000100000000000000 ; 
		block_ram[251] = 24'b010000000100000000000001 ; 
		block_ram[252] = 24'b000001100000010000010000 ; 
		block_ram[253] = 24'b001000000010000010000000 ; 
		block_ram[254] = 24'b010000000100000000000100 ; 
		block_ram[255] = 24'b000000000001011100000000 ; 
		block_ram[256] = 24'b000000000000000100000000 ; 
		block_ram[257] = 24'b000000000000000100000001 ; 
		block_ram[258] = 24'b000000000000000100000010 ; 
		block_ram[259] = 24'b000000000000000100000011 ; 
		block_ram[260] = 24'b000000000000000100000100 ; 
		block_ram[261] = 24'b000000000000000100000101 ; 
		block_ram[262] = 24'b000000000000000100000110 ; 
		block_ram[263] = 24'b000000000000000100000111 ; 
		block_ram[264] = 24'b000000000000000100001000 ; 
		block_ram[265] = 24'b000000000000000100001001 ; 
		block_ram[266] = 24'b000000000000000100001010 ; 
		block_ram[267] = 24'b000000000000000100001011 ; 
		block_ram[268] = 24'b000000000000000100001100 ; 
		block_ram[269] = 24'b000000000000000100001101 ; 
		block_ram[270] = 24'b000000000000000100001110 ; 
		block_ram[271] = 24'b001001000000010000000000 ; 
		block_ram[272] = 24'b000000000000000100010000 ; 
		block_ram[273] = 24'b000000000000000100010001 ; 
		block_ram[274] = 24'b000000000000000100010010 ; 
		block_ram[275] = 24'b000000000000000100010011 ; 
		block_ram[276] = 24'b000000000000000100010100 ; 
		block_ram[277] = 24'b000000000000000100010101 ; 
		block_ram[278] = 24'b000000000000000100010110 ; 
		block_ram[279] = 24'b000100000100000001000000 ; 
		block_ram[280] = 24'b000000000000000100011000 ; 
		block_ram[281] = 24'b000000000000000100011001 ; 
		block_ram[282] = 24'b000000000000000100011010 ; 
		block_ram[283] = 24'b000000011000000000100000 ; 
		block_ram[284] = 24'b000000000000000100011100 ; 
		block_ram[285] = 24'b100000000001100000000000 ; 
		block_ram[286] = 24'b000000100010000010000000 ; 
		block_ram[287] = 24'b000000011000000000100100 ; 
		block_ram[288] = 24'b000000000000000100100000 ; 
		block_ram[289] = 24'b000000000000000100100001 ; 
		block_ram[290] = 24'b000000000000000100100010 ; 
		block_ram[291] = 24'b000000000000000100100011 ; 
		block_ram[292] = 24'b000000000000000100100100 ; 
		block_ram[293] = 24'b000000000000000100100101 ; 
		block_ram[294] = 24'b000000000000000100100110 ; 
		block_ram[295] = 24'b100000000010001000000000 ; 
		block_ram[296] = 24'b000000000000000100101000 ; 
		block_ram[297] = 24'b000000000000000100101001 ; 
		block_ram[298] = 24'b000000000000000100101010 ; 
		block_ram[299] = 24'b000000011000000000010000 ; 
		block_ram[300] = 24'b000000000000000100101100 ; 
		block_ram[301] = 24'b010100000000000010000000 ; 
		block_ram[302] = 24'b000010000000100001000000 ; 
		block_ram[303] = 24'b000000011000000000010100 ; 
		block_ram[304] = 24'b000000000000000100110000 ; 
		block_ram[305] = 24'b000000000000000100110001 ; 
		block_ram[306] = 24'b000000000000000100110010 ; 
		block_ram[307] = 24'b000000011000000000001000 ; 
		block_ram[308] = 24'b000000000000000100110100 ; 
		block_ram[309] = 24'b000010100000010000000000 ; 
		block_ram[310] = 24'b011000000001000000000000 ; 
		block_ram[311] = 24'b000000011000000000001100 ; 
		block_ram[312] = 24'b000000000000000100111000 ; 
		block_ram[313] = 24'b000000011000000000000010 ; 
		block_ram[314] = 24'b000000011000000000000001 ; 
		block_ram[315] = 24'b000000011000000000000000 ; 
		block_ram[316] = 24'b000001000100001000000000 ; 
		block_ram[317] = 24'b000000011000000000000110 ; 
		block_ram[318] = 24'b000000011000000000000101 ; 
		block_ram[319] = 24'b000000011000000000000100 ; 
		block_ram[320] = 24'b000000000000000101000000 ; 
		block_ram[321] = 24'b000000000000000101000001 ; 
		block_ram[322] = 24'b000000000000000101000010 ; 
		block_ram[323] = 24'b000000000000000101000011 ; 
		block_ram[324] = 24'b000000000000000101000100 ; 
		block_ram[325] = 24'b000000000000000101000101 ; 
		block_ram[326] = 24'b000000000000000101000110 ; 
		block_ram[327] = 24'b000100000100000000010000 ; 
		block_ram[328] = 24'b000000000000000101001000 ; 
		block_ram[329] = 24'b000000000000000101001001 ; 
		block_ram[330] = 24'b000000000000000101001010 ; 
		block_ram[331] = 24'b010000000011000000000000 ; 
		block_ram[332] = 24'b000000000000000101001100 ; 
		block_ram[333] = 24'b000000101000001000000000 ; 
		block_ram[334] = 24'b000010000000100000100000 ; 
		block_ram[335] = 24'b000000101000001000000010 ; 
		block_ram[336] = 24'b000000000000000101010000 ; 
		block_ram[337] = 24'b000000000000000101010001 ; 
		block_ram[338] = 24'b000000000000000101010010 ; 
		block_ram[339] = 24'b000100000100000000000100 ; 
		block_ram[340] = 24'b000000000000000101010100 ; 
		block_ram[341] = 24'b000100000100000000000010 ; 
		block_ram[342] = 24'b000100000100000000000001 ; 
		block_ram[343] = 24'b000100000100000000000000 ; 
		block_ram[344] = 24'b000000000000000101011000 ; 
		block_ram[345] = 24'b000011000000000010000000 ; 
		block_ram[346] = 24'b101000000000001000000000 ; 
		block_ram[347] = 24'b000000011000000001100000 ; 
		block_ram[348] = 24'b010000010000010000000000 ; 
		block_ram[349] = 24'b000000101000001000010000 ; 
		block_ram[350] = 24'b000000100010000011000000 ; 
		block_ram[351] = 24'b000100000100000000001000 ; 
		block_ram[352] = 24'b000000000000000101100000 ; 
		block_ram[353] = 24'b000000000000000101100001 ; 
		block_ram[354] = 24'b000000000000000101100010 ; 
		block_ram[355] = 24'b001000100000000010000000 ; 
		block_ram[356] = 24'b000000000000000101100100 ; 
		block_ram[357] = 24'b000001010001000000000000 ; 
		block_ram[358] = 24'b000010000000100000001000 ; 
		block_ram[359] = 24'b000001010001000000000010 ; 
		block_ram[360] = 24'b000000000000000101101000 ; 
		block_ram[361] = 24'b100000000100010000000000 ; 
		block_ram[362] = 24'b000010000000100000000100 ; 
		block_ram[363] = 24'b000000011000000001010000 ; 
		block_ram[364] = 24'b000010000000100000000010 ; 
		block_ram[365] = 24'b000000101000001000100000 ; 
		block_ram[366] = 24'b000010000000100000000000 ; 
		block_ram[367] = 24'b000010000000100000000001 ; 
		block_ram[368] = 24'b000000000000000101110000 ; 
		block_ram[369] = 24'b010000000000101000000000 ; 
		block_ram[370] = 24'b000001000010010000000000 ; 
		block_ram[371] = 24'b000000011000000001001000 ; 
		block_ram[372] = 24'b100000001000000010000000 ; 
		block_ram[373] = 24'b000001010001000000010000 ; 
		block_ram[374] = 24'b000000110000001100000000 ; 
		block_ram[375] = 24'b000100000100000000100000 ; 
		block_ram[376] = 24'b000100100001000000000000 ; 
		block_ram[377] = 24'b000000011000000001000010 ; 
		block_ram[378] = 24'b000000011000000001000001 ; 
		block_ram[379] = 24'b000000011000000001000000 ; 
		block_ram[380] = 24'b000001000100001001000000 ; 
		block_ram[381] = 24'b001000000010000100000000 ; 
		block_ram[382] = 24'b000010000000100000010000 ; 
		block_ram[383] = 24'b000000000001011010000000 ; 
		block_ram[384] = 24'b000000000000000110000000 ; 
		block_ram[385] = 24'b000000000000000110000001 ; 
		block_ram[386] = 24'b000000000000000110000010 ; 
		block_ram[387] = 24'b000000000000000110000011 ; 
		block_ram[388] = 24'b000000000000000110000100 ; 
		block_ram[389] = 24'b000000000000000110000101 ; 
		block_ram[390] = 24'b000000000000000110000110 ; 
		block_ram[391] = 24'b000010001001000000000000 ; 
		block_ram[392] = 24'b000000000000000110001000 ; 
		block_ram[393] = 24'b000000000000000110001001 ; 
		block_ram[394] = 24'b000000000000000110001010 ; 
		block_ram[395] = 24'b000000000100101000000000 ; 
		block_ram[396] = 24'b000000000000000110001100 ; 
		block_ram[397] = 24'b010100000000000000100000 ; 
		block_ram[398] = 24'b000000100010000000010000 ; 
		block_ram[399] = 24'b000000000100101000000100 ; 
		block_ram[400] = 24'b000000000000000110010000 ; 
		block_ram[401] = 24'b000000000000000110010001 ; 
		block_ram[402] = 24'b000000000000000110010010 ; 
		block_ram[403] = 24'b110000000000010000000000 ; 
		block_ram[404] = 24'b000000000000000110010100 ; 
		block_ram[405] = 24'b001000010000001000000000 ; 
		block_ram[406] = 24'b000000100010000000001000 ; 
		block_ram[407] = 24'b000000100010000000001001 ; 
		block_ram[408] = 24'b000000000000000110011000 ; 
		block_ram[409] = 24'b000011000000000001000000 ; 
		block_ram[410] = 24'b000000100010000000000100 ; 
		block_ram[411] = 24'b000000000100101000010000 ; 
		block_ram[412] = 24'b000000100010000000000010 ; 
		block_ram[413] = 24'b000000001100010100000000 ; 
		block_ram[414] = 24'b000000100010000000000000 ; 
		block_ram[415] = 24'b000000100010000000000001 ; 
		block_ram[416] = 24'b000000000000000110100000 ; 
		block_ram[417] = 24'b000000000000000110100001 ; 
		block_ram[418] = 24'b000000000000000110100010 ; 
		block_ram[419] = 24'b001000100000000001000000 ; 
		block_ram[420] = 24'b000000000000000110100100 ; 
		block_ram[421] = 24'b010100000000000000001000 ; 
		block_ram[422] = 24'b000000010100010000000000 ; 
		block_ram[423] = 24'b000000010100010000000001 ; 
		block_ram[424] = 24'b000000000000000110101000 ; 
		block_ram[425] = 24'b010100000000000000000100 ; 
		block_ram[426] = 24'b100001000001000000000000 ; 
		block_ram[427] = 24'b000000000100101000100000 ; 
		block_ram[428] = 24'b010100000000000000000001 ; 
		block_ram[429] = 24'b010100000000000000000000 ; 
		block_ram[430] = 24'b000000010100010000001000 ; 
		block_ram[431] = 24'b010100000000000000000010 ; 
		block_ram[432] = 24'b000000000000000110110000 ; 
		block_ram[433] = 24'b000000000111000000000000 ; 
		block_ram[434] = 24'b000110000000001000000000 ; 
		block_ram[435] = 24'b000000000111000000000010 ; 
		block_ram[436] = 24'b100000001000000001000000 ; 
		block_ram[437] = 24'b000000000111000000000100 ; 
		block_ram[438] = 24'b000000010100010000010000 ; 
		block_ram[439] = 24'b000001000000100100000000 ; 
		block_ram[440] = 24'b001000000000110000000000 ; 
		block_ram[441] = 24'b000000000111000000001000 ; 
		block_ram[442] = 24'b000000011000000010000001 ; 
		block_ram[443] = 24'b000000011000000010000000 ; 
		block_ram[444] = 24'b000000100010000000100010 ; 
		block_ram[445] = 24'b010100000000000000010000 ; 
		block_ram[446] = 24'b000000100010000000100000 ; 
		block_ram[447] = 24'b000000000001011001000000 ; 
		block_ram[448] = 24'b000000000000000111000000 ; 
		block_ram[449] = 24'b000000000000000111000001 ; 
		block_ram[450] = 24'b000000000000000111000010 ; 
		block_ram[451] = 24'b001000100000000000100000 ; 
		block_ram[452] = 24'b000000000000000111000100 ; 
		block_ram[453] = 24'b000000000010110000000000 ; 
		block_ram[454] = 24'b010001000000001000000000 ; 
		block_ram[455] = 24'b000000000010110000000010 ; 
		block_ram[456] = 24'b000000000000000111001000 ; 
		block_ram[457] = 24'b000011000000000000010000 ; 
		block_ram[458] = 24'b000100001000010000000000 ; 
		block_ram[459] = 24'b000000000100101001000000 ; 
		block_ram[460] = 24'b001000000101000000000000 ; 
		block_ram[461] = 24'b000000000010110000001000 ; 
		block_ram[462] = 24'b000000100010000001010000 ; 
		block_ram[463] = 24'b100000010000000100000000 ; 
		block_ram[464] = 24'b000000000000000111010000 ; 
		block_ram[465] = 24'b000011000000000000001000 ; 
		block_ram[466] = 24'b000000010001100000000000 ; 
		block_ram[467] = 24'b000000001010001100000000 ; 
		block_ram[468] = 24'b100000001000000000100000 ; 
		block_ram[469] = 24'b000000000010110000010000 ; 
		block_ram[470] = 24'b000000010001100000000100 ; 
		block_ram[471] = 24'b000100000100000010000000 ; 
		block_ram[472] = 24'b000011000000000000000001 ; 
		block_ram[473] = 24'b000011000000000000000000 ; 
		block_ram[474] = 24'b000000010001100000001000 ; 
		block_ram[475] = 24'b000011000000000000000010 ; 
		block_ram[476] = 24'b000000100010000001000010 ; 
		block_ram[477] = 24'b000011000000000000000100 ; 
		block_ram[478] = 24'b000000100010000001000000 ; 
		block_ram[479] = 24'b000000000001011000100000 ; 
		block_ram[480] = 24'b000000000000000111100000 ; 
		block_ram[481] = 24'b001000100000000000000010 ; 
		block_ram[482] = 24'b001000100000000000000001 ; 
		block_ram[483] = 24'b001000100000000000000000 ; 
		block_ram[484] = 24'b100000001000000000010000 ; 
		block_ram[485] = 24'b000000000010110000100000 ; 
		block_ram[486] = 24'b000000010100010001000000 ; 
		block_ram[487] = 24'b001000100000000000000100 ; 
		block_ram[488] = 24'b000000010010001000000000 ; 
		block_ram[489] = 24'b000000001001100100000000 ; 
		block_ram[490] = 24'b000000010010001000000010 ; 
		block_ram[491] = 24'b001000100000000000001000 ; 
		block_ram[492] = 24'b000000010010001000000100 ; 
		block_ram[493] = 24'b010100000000000001000000 ; 
		block_ram[494] = 24'b000010000000100010000000 ; 
		block_ram[495] = 24'b000000000001011000010000 ; 
		block_ram[496] = 24'b100000001000000000000100 ; 
		block_ram[497] = 24'b000000000111000001000000 ; 
		block_ram[498] = 24'b000000010001100000100000 ; 
		block_ram[499] = 24'b001000100000000000010000 ; 
		block_ram[500] = 24'b100000001000000000000000 ; 
		block_ram[501] = 24'b100000001000000000000001 ; 
		block_ram[502] = 24'b100000001000000000000010 ; 
		block_ram[503] = 24'b000000000001011000001000 ; 
		block_ram[504] = 24'b000000010010001000010000 ; 
		block_ram[505] = 24'b000011000000000000100000 ; 
		block_ram[506] = 24'b010000000100000100000000 ; 
		block_ram[507] = 24'b000000000001011000000100 ; 
		block_ram[508] = 24'b100000001000000000001000 ; 
		block_ram[509] = 24'b000000000001011000000010 ; 
		block_ram[510] = 24'b000000000001011000000001 ; 
		block_ram[511] = 24'b000000000001011000000000 ; 
		block_ram[512] = 24'b000000000000001000000000 ; 
		block_ram[513] = 24'b000000000000001000000001 ; 
		block_ram[514] = 24'b000000000000001000000010 ; 
		block_ram[515] = 24'b000000000000001000000011 ; 
		block_ram[516] = 24'b000000000000001000000100 ; 
		block_ram[517] = 24'b000000000000001000000101 ; 
		block_ram[518] = 24'b000000000000001000000110 ; 
		block_ram[519] = 24'b000000000000001000000111 ; 
		block_ram[520] = 24'b000000000000001000001000 ; 
		block_ram[521] = 24'b000000000000001000001001 ; 
		block_ram[522] = 24'b000000000000001000001010 ; 
		block_ram[523] = 24'b000000000000001000001011 ; 
		block_ram[524] = 24'b000000000000001000001100 ; 
		block_ram[525] = 24'b000000000000001000001101 ; 
		block_ram[526] = 24'b000000000000001000001110 ; 
		block_ram[527] = 24'b010010000000000000010000 ; 
		block_ram[528] = 24'b000000000000001000010000 ; 
		block_ram[529] = 24'b000000000000001000010001 ; 
		block_ram[530] = 24'b000000000000001000010010 ; 
		block_ram[531] = 24'b000000000000001000010011 ; 
		block_ram[532] = 24'b000000000000001000010100 ; 
		block_ram[533] = 24'b000000000000001000010101 ; 
		block_ram[534] = 24'b000000000000001000010110 ; 
		block_ram[535] = 24'b010010000000000000001000 ; 
		block_ram[536] = 24'b000000000000001000011000 ; 
		block_ram[537] = 24'b000000000000001000011001 ; 
		block_ram[538] = 24'b000000000000001000011010 ; 
		block_ram[539] = 24'b010010000000000000000100 ; 
		block_ram[540] = 24'b000000000000001000011100 ; 
		block_ram[541] = 24'b010010000000000000000010 ; 
		block_ram[542] = 24'b010010000000000000000001 ; 
		block_ram[543] = 24'b010010000000000000000000 ; 
		block_ram[544] = 24'b000000000000001000100000 ; 
		block_ram[545] = 24'b000000000000001000100001 ; 
		block_ram[546] = 24'b000000000000001000100010 ; 
		block_ram[547] = 24'b000000000000001000100011 ; 
		block_ram[548] = 24'b000000000000001000100100 ; 
		block_ram[549] = 24'b000000000000001000100101 ; 
		block_ram[550] = 24'b000000000000001000100110 ; 
		block_ram[551] = 24'b100000000010000100000000 ; 
		block_ram[552] = 24'b000000000000001000101000 ; 
		block_ram[553] = 24'b000000000000001000101001 ; 
		block_ram[554] = 24'b000000000000001000101010 ; 
		block_ram[555] = 24'b000101000000000001000000 ; 
		block_ram[556] = 24'b000000000000001000101100 ; 
		block_ram[557] = 24'b000000010000110000000000 ; 
		block_ram[558] = 24'b001000001000000010000000 ; 
		block_ram[559] = 24'b000000010000110000000010 ; 
		block_ram[560] = 24'b000000000000001000110000 ; 
		block_ram[561] = 24'b000000000000001000110001 ; 
		block_ram[562] = 24'b000000000000001000110010 ; 
		block_ram[563] = 24'b001000000100010000000000 ; 
		block_ram[564] = 24'b000000000000001000110100 ; 
		block_ram[565] = 24'b000100001001000000000000 ; 
		block_ram[566] = 24'b000000110000000001000000 ; 
		block_ram[567] = 24'b000000110000000001000001 ; 
		block_ram[568] = 24'b000000000000001000111000 ; 
		block_ram[569] = 24'b100000100000000010000000 ; 
		block_ram[570] = 24'b000000000011100000000000 ; 
		block_ram[571] = 24'b000000000011100000000001 ; 
		block_ram[572] = 24'b000001000100000100000000 ; 
		block_ram[573] = 24'b000000010000110000010000 ; 
		block_ram[574] = 24'b000000000011100000000100 ; 
		block_ram[575] = 24'b010010000000000000100000 ; 
		block_ram[576] = 24'b000000000000001001000000 ; 
		block_ram[577] = 24'b000000000000001001000001 ; 
		block_ram[578] = 24'b000000000000001001000010 ; 
		block_ram[579] = 24'b000000000000001001000011 ; 
		block_ram[580] = 24'b000000000000001001000100 ; 
		block_ram[581] = 24'b000000000000001001000101 ; 
		block_ram[582] = 24'b000000000000001001000110 ; 
		block_ram[583] = 24'b001000000001100000000000 ; 
		block_ram[584] = 24'b000000000000001001001000 ; 
		block_ram[585] = 24'b000000000000001001001001 ; 
		block_ram[586] = 24'b000000000000001001001010 ; 
		block_ram[587] = 24'b000101000000000000100000 ; 
		block_ram[588] = 24'b000000000000001001001100 ; 
		block_ram[589] = 24'b000000101000000100000000 ; 
		block_ram[590] = 24'b000000000110010000000000 ; 
		block_ram[591] = 24'b000000000110010000000001 ; 
		block_ram[592] = 24'b000000000000001001010000 ; 
		block_ram[593] = 24'b000000000000001001010001 ; 
		block_ram[594] = 24'b000000000000001001010010 ; 
		block_ram[595] = 24'b000000001010000010000000 ; 
		block_ram[596] = 24'b000000000000001001010100 ; 
		block_ram[597] = 24'b100001000000010000000000 ; 
		block_ram[598] = 24'b000000110000000000100000 ; 
		block_ram[599] = 24'b000000001010000010000100 ; 
		block_ram[600] = 24'b000000000000001001011000 ; 
		block_ram[601] = 24'b000000010101000000000000 ; 
		block_ram[602] = 24'b101000000000000100000000 ; 
		block_ram[603] = 24'b000000001010000010001000 ; 
		block_ram[604] = 24'b000100000000100010000000 ; 
		block_ram[605] = 24'b000000010101000000000100 ; 
		block_ram[606] = 24'b000000000110010000010000 ; 
		block_ram[607] = 24'b010010000000000001000000 ; 
		block_ram[608] = 24'b000000000000001001100000 ; 
		block_ram[609] = 24'b000000000000001001100001 ; 
		block_ram[610] = 24'b000000000000001001100010 ; 
		block_ram[611] = 24'b000101000000000000001000 ; 
		block_ram[612] = 24'b000000000000001001100100 ; 
		block_ram[613] = 24'b000010000100000010000000 ; 
		block_ram[614] = 24'b000000110000000000010000 ; 
		block_ram[615] = 24'b000000110000000000010001 ; 
		block_ram[616] = 24'b000000000000001001101000 ; 
		block_ram[617] = 24'b000101000000000000000010 ; 
		block_ram[618] = 24'b000101000000000000000001 ; 
		block_ram[619] = 24'b000101000000000000000000 ; 
		block_ram[620] = 24'b110000000001000000000000 ; 
		block_ram[621] = 24'b000000010000110001000000 ; 
		block_ram[622] = 24'b000000000110010000100000 ; 
		block_ram[623] = 24'b000101000000000000000100 ; 
		block_ram[624] = 24'b000000000000001001110000 ; 
		block_ram[625] = 24'b010000000000100100000000 ; 
		block_ram[626] = 24'b000000110000000000000100 ; 
		block_ram[627] = 24'b000000001010000010100000 ; 
		block_ram[628] = 24'b000000110000000000000010 ; 
		block_ram[629] = 24'b000000110000000000000011 ; 
		block_ram[630] = 24'b000000110000000000000000 ; 
		block_ram[631] = 24'b000000110000000000000001 ; 
		block_ram[632] = 24'b000010001000010000000000 ; 
		block_ram[633] = 24'b000000010101000000100000 ; 
		block_ram[634] = 24'b000000000011100001000000 ; 
		block_ram[635] = 24'b000101000000000000010000 ; 
		block_ram[636] = 24'b000000110000000000001010 ; 
		block_ram[637] = 24'b001000000010001000000000 ; 
		block_ram[638] = 24'b000000110000000000001000 ; 
		block_ram[639] = 24'b000000000001010110000000 ; 
		block_ram[640] = 24'b000000000000001010000000 ; 
		block_ram[641] = 24'b000000000000001010000001 ; 
		block_ram[642] = 24'b000000000000001010000010 ; 
		block_ram[643] = 24'b000000000000001010000011 ; 
		block_ram[644] = 24'b000000000000001010000100 ; 
		block_ram[645] = 24'b000000000000001010000101 ; 
		block_ram[646] = 24'b000000000000001010000110 ; 
		block_ram[647] = 24'b000100100000010000000000 ; 
		block_ram[648] = 24'b000000000000001010001000 ; 
		block_ram[649] = 24'b000000000000001010001001 ; 
		block_ram[650] = 24'b000000000000001010001010 ; 
		block_ram[651] = 24'b000000000100100100000000 ; 
		block_ram[652] = 24'b000000000000001010001100 ; 
		block_ram[653] = 24'b000001000011000000000000 ; 
		block_ram[654] = 24'b001000001000000000100000 ; 
		block_ram[655] = 24'b000000000100100100000100 ; 
		block_ram[656] = 24'b000000000000001010010000 ; 
		block_ram[657] = 24'b000000000000001010010001 ; 
		block_ram[658] = 24'b000000000000001010010010 ; 
		block_ram[659] = 24'b000000001010000001000000 ; 
		block_ram[660] = 24'b000000000000001010010100 ; 
		block_ram[661] = 24'b001000010000000100000000 ; 
		block_ram[662] = 24'b100000000101000000000000 ; 
		block_ram[663] = 24'b000000001010000001000100 ; 
		block_ram[664] = 24'b000000000000001010011000 ; 
		block_ram[665] = 24'b100000100000000000100000 ; 
		block_ram[666] = 24'b000001010000010000000000 ; 
		block_ram[667] = 24'b000000000100100100010000 ; 
		block_ram[668] = 24'b000100000000100001000000 ; 
		block_ram[669] = 24'b000000001100011000000000 ; 
		block_ram[670] = 24'b000000100010001100000000 ; 
		block_ram[671] = 24'b010010000000000010000000 ; 
		block_ram[672] = 24'b000000000000001010100000 ; 
		block_ram[673] = 24'b000000000000001010100001 ; 
		block_ram[674] = 24'b000000000000001010100010 ; 
		block_ram[675] = 24'b010000010001000000000000 ; 
		block_ram[676] = 24'b000000000000001010100100 ; 
		block_ram[677] = 24'b000010000100000001000000 ; 
		block_ram[678] = 24'b001000001000000000001000 ; 
		block_ram[679] = 24'b000001000000101000010000 ; 
		block_ram[680] = 24'b000000000000001010101000 ; 
		block_ram[681] = 24'b100000100000000000010000 ; 
		block_ram[682] = 24'b001000001000000000000100 ; 
		block_ram[683] = 24'b000000000100100100100000 ; 
		block_ram[684] = 24'b001000001000000000000010 ; 
		block_ram[685] = 24'b000000010000110010000000 ; 
		block_ram[686] = 24'b001000001000000000000000 ; 
		block_ram[687] = 24'b001000001000000000000001 ; 
		block_ram[688] = 24'b000000000000001010110000 ; 
		block_ram[689] = 24'b100000100000000000001000 ; 
		block_ram[690] = 24'b000110000000000100000000 ; 
		block_ram[691] = 24'b000000001010000001100000 ; 
		block_ram[692] = 24'b010000000010010000000000 ; 
		block_ram[693] = 24'b000001000000101000000010 ; 
		block_ram[694] = 24'b000000110000000011000000 ; 
		block_ram[695] = 24'b000001000000101000000000 ; 
		block_ram[696] = 24'b100000100000000000000001 ; 
		block_ram[697] = 24'b100000100000000000000000 ; 
		block_ram[698] = 24'b000000000011100010000000 ; 
		block_ram[699] = 24'b100000100000000000000010 ; 
		block_ram[700] = 24'b000001000100000110000000 ; 
		block_ram[701] = 24'b100000100000000000000100 ; 
		block_ram[702] = 24'b001000001000000000010000 ; 
		block_ram[703] = 24'b000000000001010101000000 ; 
		block_ram[704] = 24'b000000000000001011000000 ; 
		block_ram[705] = 24'b000000000000001011000001 ; 
		block_ram[706] = 24'b000000000000001011000010 ; 
		block_ram[707] = 24'b000000001010000000010000 ; 
		block_ram[708] = 24'b000000000000001011000100 ; 
		block_ram[709] = 24'b000010000100000000100000 ; 
		block_ram[710] = 24'b010001000000000100000000 ; 
		block_ram[711] = 24'b000000001010000000010100 ; 
		block_ram[712] = 24'b000000000000001011001000 ; 
		block_ram[713] = 24'b011000000000010000000000 ; 
		block_ram[714] = 24'b000010100001000000000000 ; 
		block_ram[715] = 24'b000000000100100101000000 ; 
		block_ram[716] = 24'b000100000000100000010000 ; 
		block_ram[717] = 24'b000000101000000110000000 ; 
		block_ram[718] = 24'b000000000110010010000000 ; 
		block_ram[719] = 24'b100000010000001000000000 ; 
		block_ram[720] = 24'b000000000000001011010000 ; 
		block_ram[721] = 24'b000000001010000000000010 ; 
		block_ram[722] = 24'b000000001010000000000001 ; 
		block_ram[723] = 24'b000000001010000000000000 ; 
		block_ram[724] = 24'b000100000000100000001000 ; 
		block_ram[725] = 24'b000000001010000000000110 ; 
		block_ram[726] = 24'b000000001010000000000101 ; 
		block_ram[727] = 24'b000000001010000000000100 ; 
		block_ram[728] = 24'b000100000000100000000100 ; 
		block_ram[729] = 24'b000000001010000000001010 ; 
		block_ram[730] = 24'b000000001010000000001001 ; 
		block_ram[731] = 24'b000000001010000000001000 ; 
		block_ram[732] = 24'b000100000000100000000000 ; 
		block_ram[733] = 24'b000100000000100000000001 ; 
		block_ram[734] = 24'b000100000000100000000010 ; 
		block_ram[735] = 24'b000000000001010100100000 ; 
		block_ram[736] = 24'b000000000000001011100000 ; 
		block_ram[737] = 24'b000010000100000000000100 ; 
		block_ram[738] = 24'b100000000000110000000000 ; 
		block_ram[739] = 24'b000000001010000000110000 ; 
		block_ram[740] = 24'b000010000100000000000001 ; 
		block_ram[741] = 24'b000010000100000000000000 ; 
		block_ram[742] = 24'b000000110000000010010000 ; 
		block_ram[743] = 24'b000010000100000000000010 ; 
		block_ram[744] = 24'b000000010010000100000000 ; 
		block_ram[745] = 24'b000000001001101000000000 ; 
		block_ram[746] = 24'b000000010010000100000010 ; 
		block_ram[747] = 24'b000101000000000010000000 ; 
		block_ram[748] = 24'b000000010010000100000100 ; 
		block_ram[749] = 24'b000010000100000000001000 ; 
		block_ram[750] = 24'b001000001000000001000000 ; 
		block_ram[751] = 24'b000000000001010100010000 ; 
		block_ram[752] = 24'b001001000001000000000000 ; 
		block_ram[753] = 24'b000000001010000000100010 ; 
		block_ram[754] = 24'b000000001010000000100001 ; 
		block_ram[755] = 24'b000000001010000000100000 ; 
		block_ram[756] = 24'b000000110000000010000010 ; 
		block_ram[757] = 24'b000010000100000000010000 ; 
		block_ram[758] = 24'b000000110000000010000000 ; 
		block_ram[759] = 24'b000000000001010100001000 ; 
		block_ram[760] = 24'b000000010010000100010000 ; 
		block_ram[761] = 24'b100000100000000001000000 ; 
		block_ram[762] = 24'b010000000100001000000000 ; 
		block_ram[763] = 24'b000000000001010100000100 ; 
		block_ram[764] = 24'b000100000000100000100000 ; 
		block_ram[765] = 24'b000000000001010100000010 ; 
		block_ram[766] = 24'b000000000001010100000001 ; 
		block_ram[767] = 24'b000000000001010100000000 ; 
		block_ram[768] = 24'b000000000000001100000000 ; 
		block_ram[769] = 24'b000000000000001100000001 ; 
		block_ram[770] = 24'b000000000000001100000010 ; 
		block_ram[771] = 24'b000000000000001100000011 ; 
		block_ram[772] = 24'b000000000000001100000100 ; 
		block_ram[773] = 24'b000000000000001100000101 ; 
		block_ram[774] = 24'b000000000000001100000110 ; 
		block_ram[775] = 24'b100000000010000000100000 ; 
		block_ram[776] = 24'b000000000000001100001000 ; 
		block_ram[777] = 24'b000000000000001100001001 ; 
		block_ram[778] = 24'b000000000000001100001010 ; 
		block_ram[779] = 24'b000000000100100010000000 ; 
		block_ram[780] = 24'b000000000000001100001100 ; 
		block_ram[781] = 24'b000000101000000001000000 ; 
		block_ram[782] = 24'b000100010001000000000000 ; 
		block_ram[783] = 24'b000000000100100010000100 ; 
		block_ram[784] = 24'b000000000000001100010000 ; 
		block_ram[785] = 24'b000000000000001100010001 ; 
		block_ram[786] = 24'b000000000000001100010010 ; 
		block_ram[787] = 24'b000001100001000000000000 ; 
		block_ram[788] = 24'b000000000000001100010100 ; 
		block_ram[789] = 24'b001000010000000010000000 ; 
		block_ram[790] = 24'b000000001000110000000000 ; 
		block_ram[791] = 24'b000000001000110000000001 ; 
		block_ram[792] = 24'b000000000000001100011000 ; 
		block_ram[793] = 24'b000100000010010000000000 ; 
		block_ram[794] = 24'b101000000000000001000000 ; 
		block_ram[795] = 24'b000000000100100010010000 ; 
		block_ram[796] = 24'b000001000100000000100000 ; 
		block_ram[797] = 24'b000000101000000001010000 ; 
		block_ram[798] = 24'b000000001000110000001000 ; 
		block_ram[799] = 24'b010010000000000100000000 ; 
		block_ram[800] = 24'b000000000000001100100000 ; 
		block_ram[801] = 24'b000000000000001100100001 ; 
		block_ram[802] = 24'b000000000000001100100010 ; 
		block_ram[803] = 24'b100000000010000000000100 ; 
		block_ram[804] = 24'b000000000000001100100100 ; 
		block_ram[805] = 24'b100000000010000000000010 ; 
		block_ram[806] = 24'b100000000010000000000001 ; 
		block_ram[807] = 24'b100000000010000000000000 ; 
		block_ram[808] = 24'b000000000000001100101000 ; 
		block_ram[809] = 24'b001010000001000000000000 ; 
		block_ram[810] = 24'b010000100000010000000000 ; 
		block_ram[811] = 24'b000000000100100010100000 ; 
		block_ram[812] = 24'b000001000100000000010000 ; 
		block_ram[813] = 24'b000000010000110100000000 ; 
		block_ram[814] = 24'b000001000100000000010010 ; 
		block_ram[815] = 24'b100000000010000000001000 ; 
		block_ram[816] = 24'b000000000000001100110000 ; 
		block_ram[817] = 24'b010000000000100001000000 ; 
		block_ram[818] = 24'b000110000000000010000000 ; 
		block_ram[819] = 24'b000000011000001000001000 ; 
		block_ram[820] = 24'b000001000100000000001000 ; 
		block_ram[821] = 24'b000001000100000000001001 ; 
		block_ram[822] = 24'b000000001000110000100000 ; 
		block_ram[823] = 24'b100000000010000000010000 ; 
		block_ram[824] = 24'b000001000100000000000100 ; 
		block_ram[825] = 24'b000000011000001000000010 ; 
		block_ram[826] = 24'b000000000011100100000000 ; 
		block_ram[827] = 24'b000000011000001000000000 ; 
		block_ram[828] = 24'b000001000100000000000000 ; 
		block_ram[829] = 24'b000001000100000000000001 ; 
		block_ram[830] = 24'b000001000100000000000010 ; 
		block_ram[831] = 24'b000000000001010011000000 ; 
		block_ram[832] = 24'b000000000000001101000000 ; 
		block_ram[833] = 24'b000000000000001101000001 ; 
		block_ram[834] = 24'b000000000000001101000010 ; 
		block_ram[835] = 24'b000010010000010000000000 ; 
		block_ram[836] = 24'b000000000000001101000100 ; 
		block_ram[837] = 24'b000000101000000000001000 ; 
		block_ram[838] = 24'b010001000000000010000000 ; 
		block_ram[839] = 24'b000000101000000000001010 ; 
		block_ram[840] = 24'b000000000000001101001000 ; 
		block_ram[841] = 24'b000000101000000000000100 ; 
		block_ram[842] = 24'b101000000000000000010000 ; 
		block_ram[843] = 24'b000000000100100011000000 ; 
		block_ram[844] = 24'b000000101000000000000001 ; 
		block_ram[845] = 24'b000000101000000000000000 ; 
		block_ram[846] = 24'b000000000110010100000000 ; 
		block_ram[847] = 24'b000000101000000000000010 ; 
		block_ram[848] = 24'b000000000000001101010000 ; 
		block_ram[849] = 24'b010000000000100000100000 ; 
		block_ram[850] = 24'b101000000000000000001000 ; 
		block_ram[851] = 24'b000000001010000110000000 ; 
		block_ram[852] = 24'b000010000011000000000000 ; 
		block_ram[853] = 24'b000000101000000000011000 ; 
		block_ram[854] = 24'b000000001000110001000000 ; 
		block_ram[855] = 24'b000100000100001000000000 ; 
		block_ram[856] = 24'b101000000000000000000010 ; 
		block_ram[857] = 24'b000000010101000100000000 ; 
		block_ram[858] = 24'b101000000000000000000000 ; 
		block_ram[859] = 24'b101000000000000000000001 ; 
		block_ram[860] = 24'b000000101000000000010001 ; 
		block_ram[861] = 24'b000000101000000000010000 ; 
		block_ram[862] = 24'b101000000000000000000100 ; 
		block_ram[863] = 24'b000000000001010010100000 ; 
		block_ram[864] = 24'b000000000000001101100000 ; 
		block_ram[865] = 24'b010000000000100000010000 ; 
		block_ram[866] = 24'b000000001101000000000000 ; 
		block_ram[867] = 24'b000000001101000000000001 ; 
		block_ram[868] = 24'b001100000000010000000000 ; 
		block_ram[869] = 24'b000000101000000000101000 ; 
		block_ram[870] = 24'b000000001101000000000100 ; 
		block_ram[871] = 24'b100000000010000001000000 ; 
		block_ram[872] = 24'b000000010010000010000000 ; 
		block_ram[873] = 24'b000000010010000010000001 ; 
		block_ram[874] = 24'b000000001101000000001000 ; 
		block_ram[875] = 24'b000101000000000100000000 ; 
		block_ram[876] = 24'b000000010010000010000100 ; 
		block_ram[877] = 24'b000000101000000000100000 ; 
		block_ram[878] = 24'b000010000000101000000000 ; 
		block_ram[879] = 24'b000000000001010010010000 ; 
		block_ram[880] = 24'b010000000000100000000001 ; 
		block_ram[881] = 24'b010000000000100000000000 ; 
		block_ram[882] = 24'b000000001101000000010000 ; 
		block_ram[883] = 24'b010000000000100000000010 ; 
		block_ram[884] = 24'b000000110000000100000010 ; 
		block_ram[885] = 24'b010000000000100000000100 ; 
		block_ram[886] = 24'b000000110000000100000000 ; 
		block_ram[887] = 24'b000000000001010010001000 ; 
		block_ram[888] = 24'b000000010010000010010000 ; 
		block_ram[889] = 24'b010000000000100000001000 ; 
		block_ram[890] = 24'b101000000000000000100000 ; 
		block_ram[891] = 24'b000000000001010010000100 ; 
		block_ram[892] = 24'b000001000100000001000000 ; 
		block_ram[893] = 24'b000000000001010010000010 ; 
		block_ram[894] = 24'b000000000001010010000001 ; 
		block_ram[895] = 24'b000000000001010010000000 ; 
		block_ram[896] = 24'b000000000000001110000000 ; 
		block_ram[897] = 24'b000000000000001110000001 ; 
		block_ram[898] = 24'b000000000000001110000010 ; 
		block_ram[899] = 24'b000000000100100000001000 ; 
		block_ram[900] = 24'b000000000000001110000100 ; 
		block_ram[901] = 24'b001000010000000000010000 ; 
		block_ram[902] = 24'b010001000000000001000000 ; 
		block_ram[903] = 24'b000000000100100000001100 ; 
		block_ram[904] = 24'b000000000000001110001000 ; 
		block_ram[905] = 24'b000000000100100000000010 ; 
		block_ram[906] = 24'b000000000100100000000001 ; 
		block_ram[907] = 24'b000000000100100000000000 ; 
		block_ram[908] = 24'b100010000000010000000000 ; 
		block_ram[909] = 24'b000000000100100000000110 ; 
		block_ram[910] = 24'b000000000100100000000101 ; 
		block_ram[911] = 24'b000000000100100000000100 ; 
		block_ram[912] = 24'b000000000000001110010000 ; 
		block_ram[913] = 24'b001000010000000000000100 ; 
		block_ram[914] = 24'b000110000000000000100000 ; 
		block_ram[915] = 24'b000000000100100000011000 ; 
		block_ram[916] = 24'b001000010000000000000001 ; 
		block_ram[917] = 24'b001000010000000000000000 ; 
		block_ram[918] = 24'b000000001000110010000000 ; 
		block_ram[919] = 24'b001000010000000000000010 ; 
		block_ram[920] = 24'b010000001001000000000000 ; 
		block_ram[921] = 24'b000000000100100000010010 ; 
		block_ram[922] = 24'b000000000100100000010001 ; 
		block_ram[923] = 24'b000000000100100000010000 ; 
		block_ram[924] = 24'b000000100010001000000010 ; 
		block_ram[925] = 24'b001000010000000000001000 ; 
		block_ram[926] = 24'b000000100010001000000000 ; 
		block_ram[927] = 24'b000000000001010001100000 ; 
		block_ram[928] = 24'b000000000000001110100000 ; 
		block_ram[929] = 24'b000001001000010000000000 ; 
		block_ram[930] = 24'b000110000000000000010000 ; 
		block_ram[931] = 24'b000000000100100000101000 ; 
		block_ram[932] = 24'b000000100001100000000000 ; 
		block_ram[933] = 24'b000000100001100000000001 ; 
		block_ram[934] = 24'b000000010100011000000000 ; 
		block_ram[935] = 24'b100000000010000010000000 ; 
		block_ram[936] = 24'b000000010010000001000000 ; 
		block_ram[937] = 24'b000000000100100000100010 ; 
		block_ram[938] = 24'b000000000100100000100001 ; 
		block_ram[939] = 24'b000000000100100000100000 ; 
		block_ram[940] = 24'b000000010010000001000100 ; 
		block_ram[941] = 24'b010100000000001000000000 ; 
		block_ram[942] = 24'b001000001000000100000000 ; 
		block_ram[943] = 24'b000000000001010001010000 ; 
		block_ram[944] = 24'b000110000000000000000010 ; 
		block_ram[945] = 24'b000000000111001000000000 ; 
		block_ram[946] = 24'b000110000000000000000000 ; 
		block_ram[947] = 24'b000110000000000000000001 ; 
		block_ram[948] = 24'b000000100001100000010000 ; 
		block_ram[949] = 24'b001000010000000000100000 ; 
		block_ram[950] = 24'b000110000000000000000100 ; 
		block_ram[951] = 24'b000000000001010001001000 ; 
		block_ram[952] = 24'b000000010010000001010000 ; 
		block_ram[953] = 24'b100000100000000100000000 ; 
		block_ram[954] = 24'b000110000000000000001000 ; 
		block_ram[955] = 24'b000000000001010001000100 ; 
		block_ram[956] = 24'b000001000100000010000000 ; 
		block_ram[957] = 24'b000000000001010001000010 ; 
		block_ram[958] = 24'b000000000001010001000001 ; 
		block_ram[959] = 24'b000000000001010001000000 ; 
		block_ram[960] = 24'b000000000000001111000000 ; 
		block_ram[961] = 24'b100100000001000000000000 ; 
		block_ram[962] = 24'b010001000000000000000100 ; 
		block_ram[963] = 24'b000000000100100001001000 ; 
		block_ram[964] = 24'b010001000000000000000010 ; 
		block_ram[965] = 24'b000000000010111000000000 ; 
		block_ram[966] = 24'b010001000000000000000000 ; 
		block_ram[967] = 24'b010001000000000000000001 ; 
		block_ram[968] = 24'b000000010010000000100000 ; 
		block_ram[969] = 24'b000000000100100001000010 ; 
		block_ram[970] = 24'b000000000100100001000001 ; 
		block_ram[971] = 24'b000000000100100001000000 ; 
		block_ram[972] = 24'b000000010010000000100100 ; 
		block_ram[973] = 24'b000000101000000010000000 ; 
		block_ram[974] = 24'b010001000000000000001000 ; 
		block_ram[975] = 24'b000000000001010000110000 ; 
		block_ram[976] = 24'b000000100100010000000000 ; 
		block_ram[977] = 24'b000000001010000100000010 ; 
		block_ram[978] = 24'b000000001010000100000001 ; 
		block_ram[979] = 24'b000000001010000100000000 ; 
		block_ram[980] = 24'b000000100100010000000100 ; 
		block_ram[981] = 24'b001000010000000001000000 ; 
		block_ram[982] = 24'b010001000000000000010000 ; 
		block_ram[983] = 24'b000000000001010000101000 ; 
		block_ram[984] = 24'b000000010010000000110000 ; 
		block_ram[985] = 24'b000011000000001000000000 ; 
		block_ram[986] = 24'b101000000000000010000000 ; 
		block_ram[987] = 24'b000000000001010000100100 ; 
		block_ram[988] = 24'b000100000000100100000000 ; 
		block_ram[989] = 24'b000000000001010000100010 ; 
		block_ram[990] = 24'b000000000001010000100001 ; 
		block_ram[991] = 24'b000000000001010000100000 ; 
		block_ram[992] = 24'b000000010010000000001000 ; 
		block_ram[993] = 24'b000000010010000000001001 ; 
		block_ram[994] = 24'b000000001101000010000000 ; 
		block_ram[995] = 24'b001000100000001000000000 ; 
		block_ram[996] = 24'b000000010010000000001100 ; 
		block_ram[997] = 24'b000010000100000100000000 ; 
		block_ram[998] = 24'b010001000000000000100000 ; 
		block_ram[999] = 24'b000000000001010000011000 ; 
		block_ram[1000] = 24'b000000010010000000000000 ; 
		block_ram[1001] = 24'b000000010010000000000001 ; 
		block_ram[1002] = 24'b000000010010000000000010 ; 
		block_ram[1003] = 24'b000000000001010000010100 ; 
		block_ram[1004] = 24'b000000010010000000000100 ; 
		block_ram[1005] = 24'b000000000001010000010010 ; 
		block_ram[1006] = 24'b000000000001010000010001 ; 
		block_ram[1007] = 24'b000000000001010000010000 ; 
		block_ram[1008] = 24'b000000010010000000011000 ; 
		block_ram[1009] = 24'b010000000000100010000000 ; 
		block_ram[1010] = 24'b000110000000000001000000 ; 
		block_ram[1011] = 24'b000000000001010000001100 ; 
		block_ram[1012] = 24'b100000001000001000000000 ; 
		block_ram[1013] = 24'b000000000001010000001010 ; 
		block_ram[1014] = 24'b000000000001010000001001 ; 
		block_ram[1015] = 24'b000000000001010000001000 ; 
		block_ram[1016] = 24'b000000010010000000010000 ; 
		block_ram[1017] = 24'b000000000001010000000110 ; 
		block_ram[1018] = 24'b000000000001010000000101 ; 
		block_ram[1019] = 24'b000000000001010000000100 ; 
		block_ram[1020] = 24'b000000000001010000000011 ; 
		block_ram[1021] = 24'b000000000001010000000010 ; 
		block_ram[1022] = 24'b000000000001010000000001 ; 
		block_ram[1023] = 24'b000000000001010000000000 ; 
		block_ram[1024] = 24'b000000000000010000000000 ; 
		block_ram[1025] = 24'b000000000000010000000001 ; 
		block_ram[1026] = 24'b000000000000010000000010 ; 
		block_ram[1027] = 24'b000000000000010000000011 ; 
		block_ram[1028] = 24'b000000000000010000000100 ; 
		block_ram[1029] = 24'b000000000000010000000101 ; 
		block_ram[1030] = 24'b000000000000010000000110 ; 
		block_ram[1031] = 24'b000000000000010000000111 ; 
		block_ram[1032] = 24'b000000000000010000001000 ; 
		block_ram[1033] = 24'b000000000000010000001001 ; 
		block_ram[1034] = 24'b000000000000010000001010 ; 
		block_ram[1035] = 24'b000000000000010000001011 ; 
		block_ram[1036] = 24'b000000000000010000001100 ; 
		block_ram[1037] = 24'b000000000000010000001101 ; 
		block_ram[1038] = 24'b000000000000010000001110 ; 
		block_ram[1039] = 24'b001001000000000100000000 ; 
		block_ram[1040] = 24'b000000000000010000010000 ; 
		block_ram[1041] = 24'b000000000000010000010001 ; 
		block_ram[1042] = 24'b000000000000010000010010 ; 
		block_ram[1043] = 24'b000000000000010000010011 ; 
		block_ram[1044] = 24'b000000000000010000010100 ; 
		block_ram[1045] = 24'b000000000000010000010101 ; 
		block_ram[1046] = 24'b000000000000010000010110 ; 
		block_ram[1047] = 24'b000000010011000000000000 ; 
		block_ram[1048] = 24'b000000000000010000011000 ; 
		block_ram[1049] = 24'b000000000000010000011001 ; 
		block_ram[1050] = 24'b000000000000010000011010 ; 
		block_ram[1051] = 24'b000000100000100001000000 ; 
		block_ram[1052] = 24'b000000000000010000011100 ; 
		block_ram[1053] = 24'b000000001100000010000000 ; 
		block_ram[1054] = 24'b100100000000000000100000 ; 
		block_ram[1055] = 24'b000000001100000010000010 ; 
		block_ram[1056] = 24'b000000000000010000100000 ; 
		block_ram[1057] = 24'b000000000000010000100001 ; 
		block_ram[1058] = 24'b000000000000010000100010 ; 
		block_ram[1059] = 24'b000000000000010000100011 ; 
		block_ram[1060] = 24'b000000000000010000100100 ; 
		block_ram[1061] = 24'b000000000000010000100101 ; 
		block_ram[1062] = 24'b000000000000010000100110 ; 
		block_ram[1063] = 24'b010000001000000001000000 ; 
		block_ram[1064] = 24'b000000000000010000101000 ; 
		block_ram[1065] = 24'b000000000000010000101001 ; 
		block_ram[1066] = 24'b000000000000010000101010 ; 
		block_ram[1067] = 24'b000010000010000010000000 ; 
		block_ram[1068] = 24'b000000000000010000101100 ; 
		block_ram[1069] = 24'b000000010000101000000000 ; 
		block_ram[1070] = 24'b100100000000000000010000 ; 
		block_ram[1071] = 24'b000000010000101000000010 ; 
		block_ram[1072] = 24'b000000000000010000110000 ; 
		block_ram[1073] = 24'b000000000000010000110001 ; 
		block_ram[1074] = 24'b000000000000010000110010 ; 
		block_ram[1075] = 24'b001000000100001000000000 ; 
		block_ram[1076] = 24'b000000000000010000110100 ; 
		block_ram[1077] = 24'b000010100000000100000000 ; 
		block_ram[1078] = 24'b100100000000000000001000 ; 
		block_ram[1079] = 24'b000000010011000000100000 ; 
		block_ram[1080] = 24'b000000000000010000111000 ; 
		block_ram[1081] = 24'b010001000001000000000000 ; 
		block_ram[1082] = 24'b100100000000000000000100 ; 
		block_ram[1083] = 24'b000000011000010100000000 ; 
		block_ram[1084] = 24'b100100000000000000000010 ; 
		block_ram[1085] = 24'b000000001100000010100000 ; 
		block_ram[1086] = 24'b100100000000000000000000 ; 
		block_ram[1087] = 24'b100100000000000000000001 ; 
		block_ram[1088] = 24'b000000000000010001000000 ; 
		block_ram[1089] = 24'b000000000000010001000001 ; 
		block_ram[1090] = 24'b000000000000010001000010 ; 
		block_ram[1091] = 24'b000000000000010001000011 ; 
		block_ram[1092] = 24'b000000000000010001000100 ; 
		block_ram[1093] = 24'b000000000000010001000101 ; 
		block_ram[1094] = 24'b000000000000010001000110 ; 
		block_ram[1095] = 24'b010000001000000000100000 ; 
		block_ram[1096] = 24'b000000000000010001001000 ; 
		block_ram[1097] = 24'b000000000000010001001001 ; 
		block_ram[1098] = 24'b000000000000010001001010 ; 
		block_ram[1099] = 24'b000000100000100000010000 ; 
		block_ram[1100] = 24'b000000000000010001001100 ; 
		block_ram[1101] = 24'b000110000001000000000000 ; 
		block_ram[1102] = 24'b000000000110001000000000 ; 
		block_ram[1103] = 24'b000000000110001000000001 ; 
		block_ram[1104] = 24'b000000000000010001010000 ; 
		block_ram[1105] = 24'b000000000000010001010001 ; 
		block_ram[1106] = 24'b000000000000010001010010 ; 
		block_ram[1107] = 24'b000000100000100000001000 ; 
		block_ram[1108] = 24'b000000000000010001010100 ; 
		block_ram[1109] = 24'b100001000000001000000000 ; 
		block_ram[1110] = 24'b001010000000000010000000 ; 
		block_ram[1111] = 24'b000000010011000001000000 ; 
		block_ram[1112] = 24'b000000000000010001011000 ; 
		block_ram[1113] = 24'b000000100000100000000010 ; 
		block_ram[1114] = 24'b000000100000100000000001 ; 
		block_ram[1115] = 24'b000000100000100000000000 ; 
		block_ram[1116] = 24'b010000010000000100000000 ; 
		block_ram[1117] = 24'b000000001100000011000000 ; 
		block_ram[1118] = 24'b000000000110001000010000 ; 
		block_ram[1119] = 24'b000000100000100000000100 ; 
		block_ram[1120] = 24'b000000000000010001100000 ; 
		block_ram[1121] = 24'b000000000000010001100001 ; 
		block_ram[1122] = 24'b000000000000010001100010 ; 
		block_ram[1123] = 24'b010000001000000000000100 ; 
		block_ram[1124] = 24'b000000000000010001100100 ; 
		block_ram[1125] = 24'b010000001000000000000010 ; 
		block_ram[1126] = 24'b010000001000000000000001 ; 
		block_ram[1127] = 24'b010000001000000000000000 ; 
		block_ram[1128] = 24'b000000000000010001101000 ; 
		block_ram[1129] = 24'b100000000100000100000000 ; 
		block_ram[1130] = 24'b001000010001000000000000 ; 
		block_ram[1131] = 24'b000000100000100000110000 ; 
		block_ram[1132] = 24'b000001100000000010000000 ; 
		block_ram[1133] = 24'b000000010000101001000000 ; 
		block_ram[1134] = 24'b000000000110001000100000 ; 
		block_ram[1135] = 24'b010000001000000000001000 ; 
		block_ram[1136] = 24'b000000000000010001110000 ; 
		block_ram[1137] = 24'b000100010000000010000000 ; 
		block_ram[1138] = 24'b000001000010000100000000 ; 
		block_ram[1139] = 24'b000000100000100000101000 ; 
		block_ram[1140] = 24'b000000000101100000000000 ; 
		block_ram[1141] = 24'b000000000101100000000001 ; 
		block_ram[1142] = 24'b000000000101100000000010 ; 
		block_ram[1143] = 24'b010000001000000000010000 ; 
		block_ram[1144] = 24'b000010001000001000000000 ; 
		block_ram[1145] = 24'b000000100000100000100010 ; 
		block_ram[1146] = 24'b000000100000100000100001 ; 
		block_ram[1147] = 24'b000000100000100000100000 ; 
		block_ram[1148] = 24'b000000000101100000001000 ; 
		block_ram[1149] = 24'b001000000010010000000000 ; 
		block_ram[1150] = 24'b100100000000000001000000 ; 
		block_ram[1151] = 24'b000000000001001110000000 ; 
		block_ram[1152] = 24'b000000000000010010000000 ; 
		block_ram[1153] = 24'b000000000000010010000001 ; 
		block_ram[1154] = 24'b000000000000010010000010 ; 
		block_ram[1155] = 24'b000000000000010010000011 ; 
		block_ram[1156] = 24'b000000000000010010000100 ; 
		block_ram[1157] = 24'b000000000000010010000101 ; 
		block_ram[1158] = 24'b000000000000010010000110 ; 
		block_ram[1159] = 24'b000100100000001000000000 ; 
		block_ram[1160] = 24'b000000000000010010001000 ; 
		block_ram[1161] = 24'b000000000000010010001001 ; 
		block_ram[1162] = 24'b000000000000010010001010 ; 
		block_ram[1163] = 24'b000010000010000000100000 ; 
		block_ram[1164] = 24'b000000000000010010001100 ; 
		block_ram[1165] = 24'b000000001100000000010000 ; 
		block_ram[1166] = 24'b010000000001100000000000 ; 
		block_ram[1167] = 24'b000000001100000000010010 ; 
		block_ram[1168] = 24'b000000000000010010010000 ; 
		block_ram[1169] = 24'b000000000000010010010001 ; 
		block_ram[1170] = 24'b000000000000010010010010 ; 
		block_ram[1171] = 24'b110000000000000100000000 ; 
		block_ram[1172] = 24'b000000000000010010010100 ; 
		block_ram[1173] = 24'b000000001100000000001000 ; 
		block_ram[1174] = 24'b001010000000000001000000 ; 
		block_ram[1175] = 24'b000000001100000000001010 ; 
		block_ram[1176] = 24'b000000000000010010011000 ; 
		block_ram[1177] = 24'b000000001100000000000100 ; 
		block_ram[1178] = 24'b000001010000001000000000 ; 
		block_ram[1179] = 24'b000000001100000000000110 ; 
		block_ram[1180] = 24'b000000001100000000000001 ; 
		block_ram[1181] = 24'b000000001100000000000000 ; 
		block_ram[1182] = 24'b000000001100000000000011 ; 
		block_ram[1183] = 24'b000000001100000000000010 ; 
		block_ram[1184] = 24'b000000000000010010100000 ; 
		block_ram[1185] = 24'b000000000000010010100001 ; 
		block_ram[1186] = 24'b000000000000010010100010 ; 
		block_ram[1187] = 24'b000010000010000000001000 ; 
		block_ram[1188] = 24'b000000000000010010100100 ; 
		block_ram[1189] = 24'b101000000001000000000000 ; 
		block_ram[1190] = 24'b000000010100000100000000 ; 
		block_ram[1191] = 24'b000000010100000100000001 ; 
		block_ram[1192] = 24'b000000000000010010101000 ; 
		block_ram[1193] = 24'b000010000010000000000010 ; 
		block_ram[1194] = 24'b000010000010000000000001 ; 
		block_ram[1195] = 24'b000010000010000000000000 ; 
		block_ram[1196] = 24'b000001100000000001000000 ; 
		block_ram[1197] = 24'b000000001100000000110000 ; 
		block_ram[1198] = 24'b000000010100000100001000 ; 
		block_ram[1199] = 24'b000010000010000000000100 ; 
		block_ram[1200] = 24'b000000000000010010110000 ; 
		block_ram[1201] = 24'b000100010000000001000000 ; 
		block_ram[1202] = 24'b000000101001000000000000 ; 
		block_ram[1203] = 24'b000000101001000000000001 ; 
		block_ram[1204] = 24'b010000000010001000000000 ; 
		block_ram[1205] = 24'b000000001100000000101000 ; 
		block_ram[1206] = 24'b000000010100000100010000 ; 
		block_ram[1207] = 24'b000001000000110000000000 ; 
		block_ram[1208] = 24'b001000000000100100000000 ; 
		block_ram[1209] = 24'b000000001100000000100100 ; 
		block_ram[1210] = 24'b000000101001000000001000 ; 
		block_ram[1211] = 24'b000010000010000000010000 ; 
		block_ram[1212] = 24'b000000001100000000100001 ; 
		block_ram[1213] = 24'b000000001100000000100000 ; 
		block_ram[1214] = 24'b100100000000000010000000 ; 
		block_ram[1215] = 24'b000000000001001101000000 ; 
		block_ram[1216] = 24'b000000000000010011000000 ; 
		block_ram[1217] = 24'b000000000000010011000001 ; 
		block_ram[1218] = 24'b000000000000010011000010 ; 
		block_ram[1219] = 24'b000001000101000000000000 ; 
		block_ram[1220] = 24'b000000000000010011000100 ; 
		block_ram[1221] = 24'b000000000010100100000000 ; 
		block_ram[1222] = 24'b001010000000000000010000 ; 
		block_ram[1223] = 24'b000000000010100100000010 ; 
		block_ram[1224] = 24'b000000000000010011001000 ; 
		block_ram[1225] = 24'b011000000000001000000000 ; 
		block_ram[1226] = 24'b000100001000000100000000 ; 
		block_ram[1227] = 24'b000000100000100010010000 ; 
		block_ram[1228] = 24'b000001100000000000100000 ; 
		block_ram[1229] = 24'b000000000010100100001000 ; 
		block_ram[1230] = 24'b000000000110001010000000 ; 
		block_ram[1231] = 24'b100000010000010000000000 ; 
		block_ram[1232] = 24'b000000000000010011010000 ; 
		block_ram[1233] = 24'b000100010000000000100000 ; 
		block_ram[1234] = 24'b001010000000000000000100 ; 
		block_ram[1235] = 24'b000000001010011000000000 ; 
		block_ram[1236] = 24'b001010000000000000000010 ; 
		block_ram[1237] = 24'b000000000010100100010000 ; 
		block_ram[1238] = 24'b001010000000000000000000 ; 
		block_ram[1239] = 24'b001010000000000000000001 ; 
		block_ram[1240] = 24'b100000000011000000000000 ; 
		block_ram[1241] = 24'b000000001100000001000100 ; 
		block_ram[1242] = 24'b000000100000100010000001 ; 
		block_ram[1243] = 24'b000000100000100010000000 ; 
		block_ram[1244] = 24'b000000001100000001000001 ; 
		block_ram[1245] = 24'b000000001100000001000000 ; 
		block_ram[1246] = 24'b001010000000000000001000 ; 
		block_ram[1247] = 24'b000000000001001100100000 ; 
		block_ram[1248] = 24'b000000000000010011100000 ; 
		block_ram[1249] = 24'b000100010000000000010000 ; 
		block_ram[1250] = 24'b100000000000101000000000 ; 
		block_ram[1251] = 24'b000001000101000000100000 ; 
		block_ram[1252] = 24'b000001100000000000001000 ; 
		block_ram[1253] = 24'b000000000010100100100000 ; 
		block_ram[1254] = 24'b000000010100000101000000 ; 
		block_ram[1255] = 24'b010000001000000010000000 ; 
		block_ram[1256] = 24'b000001100000000000000100 ; 
		block_ram[1257] = 24'b000000001001110000000000 ; 
		block_ram[1258] = 24'b000001100000000000000110 ; 
		block_ram[1259] = 24'b000010000010000001000000 ; 
		block_ram[1260] = 24'b000001100000000000000000 ; 
		block_ram[1261] = 24'b000001100000000000000001 ; 
		block_ram[1262] = 24'b000001100000000000000010 ; 
		block_ram[1263] = 24'b000000000001001100010000 ; 
		block_ram[1264] = 24'b000100010000000000000001 ; 
		block_ram[1265] = 24'b000100010000000000000000 ; 
		block_ram[1266] = 24'b000000101001000001000000 ; 
		block_ram[1267] = 24'b000100010000000000000010 ; 
		block_ram[1268] = 24'b000000000101100010000000 ; 
		block_ram[1269] = 24'b000100010000000000000100 ; 
		block_ram[1270] = 24'b001010000000000000100000 ; 
		block_ram[1271] = 24'b000000000001001100001000 ; 
		block_ram[1272] = 24'b000001100000000000010100 ; 
		block_ram[1273] = 24'b000100010000000000001000 ; 
		block_ram[1274] = 24'b010000000100010000000000 ; 
		block_ram[1275] = 24'b000000000001001100000100 ; 
		block_ram[1276] = 24'b000001100000000000010000 ; 
		block_ram[1277] = 24'b000000000001001100000010 ; 
		block_ram[1278] = 24'b000000000001001100000001 ; 
		block_ram[1279] = 24'b000000000001001100000000 ; 
		block_ram[1280] = 24'b000000000000010100000000 ; 
		block_ram[1281] = 24'b000000000000010100000001 ; 
		block_ram[1282] = 24'b000000000000010100000010 ; 
		block_ram[1283] = 24'b000000000000010100000011 ; 
		block_ram[1284] = 24'b000000000000010100000100 ; 
		block_ram[1285] = 24'b000000000000010100000101 ; 
		block_ram[1286] = 24'b000000000000010100000110 ; 
		block_ram[1287] = 24'b001001000000000000001000 ; 
		block_ram[1288] = 24'b000000000000010100001000 ; 
		block_ram[1289] = 24'b000000000000010100001001 ; 
		block_ram[1290] = 24'b000000000000010100001010 ; 
		block_ram[1291] = 24'b001001000000000000000100 ; 
		block_ram[1292] = 24'b000000000000010100001100 ; 
		block_ram[1293] = 24'b001001000000000000000010 ; 
		block_ram[1294] = 24'b001001000000000000000001 ; 
		block_ram[1295] = 24'b001001000000000000000000 ; 
		block_ram[1296] = 24'b000000000000010100010000 ; 
		block_ram[1297] = 24'b000000000000010100010001 ; 
		block_ram[1298] = 24'b000000000000010100010010 ; 
		block_ram[1299] = 24'b110000000000000010000000 ; 
		block_ram[1300] = 24'b000000000000010100010100 ; 
		block_ram[1301] = 24'b000010100000000000100000 ; 
		block_ram[1302] = 24'b000000001000101000000000 ; 
		block_ram[1303] = 24'b000000001000101000000001 ; 
		block_ram[1304] = 24'b000000000000010100011000 ; 
		block_ram[1305] = 24'b000100000010001000000000 ; 
		block_ram[1306] = 24'b000010000101000000000000 ; 
		block_ram[1307] = 24'b000000011000010000100000 ; 
		block_ram[1308] = 24'b010000010000000001000000 ; 
		block_ram[1309] = 24'b000000001100000110000000 ; 
		block_ram[1310] = 24'b000000001000101000001000 ; 
		block_ram[1311] = 24'b001001000000000000010000 ; 
		block_ram[1312] = 24'b000000000000010100100000 ; 
		block_ram[1313] = 24'b000000000000010100100001 ; 
		block_ram[1314] = 24'b000000000000010100100010 ; 
		block_ram[1315] = 24'b000100000001100000000000 ; 
		block_ram[1316] = 24'b000000000000010100100100 ; 
		block_ram[1317] = 24'b000010100000000000010000 ; 
		block_ram[1318] = 24'b000000010100000010000000 ; 
		block_ram[1319] = 24'b000000010100000010000001 ; 
		block_ram[1320] = 24'b000000000000010100101000 ; 
		block_ram[1321] = 24'b100000000100000001000000 ; 
		block_ram[1322] = 24'b010000100000001000000000 ; 
		block_ram[1323] = 24'b000000011000010000010000 ; 
		block_ram[1324] = 24'b000000001011000000000000 ; 
		block_ram[1325] = 24'b000000001011000000000001 ; 
		block_ram[1326] = 24'b000000001011000000000010 ; 
		block_ram[1327] = 24'b001001000000000000100000 ; 
		block_ram[1328] = 24'b000000000000010100110000 ; 
		block_ram[1329] = 24'b000010100000000000000100 ; 
		block_ram[1330] = 24'b000001000010000001000000 ; 
		block_ram[1331] = 24'b000000011000010000001000 ; 
		block_ram[1332] = 24'b000010100000000000000001 ; 
		block_ram[1333] = 24'b000010100000000000000000 ; 
		block_ram[1334] = 24'b000000001000101000100000 ; 
		block_ram[1335] = 24'b000010100000000000000010 ; 
		block_ram[1336] = 24'b001000000000100010000000 ; 
		block_ram[1337] = 24'b000000011000010000000010 ; 
		block_ram[1338] = 24'b000000011000010000000001 ; 
		block_ram[1339] = 24'b000000011000010000000000 ; 
		block_ram[1340] = 24'b000000001011000000010000 ; 
		block_ram[1341] = 24'b000010100000000000001000 ; 
		block_ram[1342] = 24'b100100000000000100000000 ; 
		block_ram[1343] = 24'b000000000001001011000000 ; 
		block_ram[1344] = 24'b000000000000010101000000 ; 
		block_ram[1345] = 24'b000000000000010101000001 ; 
		block_ram[1346] = 24'b000000000000010101000010 ; 
		block_ram[1347] = 24'b000010010000001000000000 ; 
		block_ram[1348] = 24'b000000000000010101000100 ; 
		block_ram[1349] = 24'b000000000010100010000000 ; 
		block_ram[1350] = 24'b100000100001000000000000 ; 
		block_ram[1351] = 24'b000000000010100010000010 ; 
		block_ram[1352] = 24'b000000000000010101001000 ; 
		block_ram[1353] = 24'b100000000100000000100000 ; 
		block_ram[1354] = 24'b000100001000000010000000 ; 
		block_ram[1355] = 24'b000000100000100100010000 ; 
		block_ram[1356] = 24'b010000010000000000010000 ; 
		block_ram[1357] = 24'b000000000010100010001000 ; 
		block_ram[1358] = 24'b000000000110001100000000 ; 
		block_ram[1359] = 24'b001001000000000001000000 ; 
		block_ram[1360] = 24'b000000000000010101010000 ; 
		block_ram[1361] = 24'b001000001001000000000000 ; 
		block_ram[1362] = 24'b000001000010000000100000 ; 
		block_ram[1363] = 24'b000000100000100100001000 ; 
		block_ram[1364] = 24'b010000010000000000001000 ; 
		block_ram[1365] = 24'b000000000010100010010000 ; 
		block_ram[1366] = 24'b000000001000101001000000 ; 
		block_ram[1367] = 24'b000100000100010000000000 ; 
		block_ram[1368] = 24'b010000010000000000000100 ; 
		block_ram[1369] = 24'b000000100000100100000010 ; 
		block_ram[1370] = 24'b000000100000100100000001 ; 
		block_ram[1371] = 24'b000000100000100100000000 ; 
		block_ram[1372] = 24'b010000010000000000000000 ; 
		block_ram[1373] = 24'b010000010000000000000001 ; 
		block_ram[1374] = 24'b010000010000000000000010 ; 
		block_ram[1375] = 24'b000000000001001010100000 ; 
		block_ram[1376] = 24'b000000000000010101100000 ; 
		block_ram[1377] = 24'b100000000100000000001000 ; 
		block_ram[1378] = 24'b000001000010000000010000 ; 
		block_ram[1379] = 24'b000001000010000000010001 ; 
		block_ram[1380] = 24'b001100000000001000000000 ; 
		block_ram[1381] = 24'b000000000010100010100000 ; 
		block_ram[1382] = 24'b000000010100000011000000 ; 
		block_ram[1383] = 24'b010000001000000100000000 ; 
		block_ram[1384] = 24'b100000000100000000000001 ; 
		block_ram[1385] = 24'b100000000100000000000000 ; 
		block_ram[1386] = 24'b000001000010000000011000 ; 
		block_ram[1387] = 24'b100000000100000000000010 ; 
		block_ram[1388] = 24'b000000001011000001000000 ; 
		block_ram[1389] = 24'b100000000100000000000100 ; 
		block_ram[1390] = 24'b000010000000110000000000 ; 
		block_ram[1391] = 24'b000000000001001010010000 ; 
		block_ram[1392] = 24'b000001000010000000000010 ; 
		block_ram[1393] = 24'b000001000010000000000011 ; 
		block_ram[1394] = 24'b000001000010000000000000 ; 
		block_ram[1395] = 24'b000001000010000000000001 ; 
		block_ram[1396] = 24'b000000000101100100000000 ; 
		block_ram[1397] = 24'b000010100000000001000000 ; 
		block_ram[1398] = 24'b000001000010000000000100 ; 
		block_ram[1399] = 24'b000000000001001010001000 ; 
		block_ram[1400] = 24'b000001000010000000001010 ; 
		block_ram[1401] = 24'b100000000100000000010000 ; 
		block_ram[1402] = 24'b000001000010000000001000 ; 
		block_ram[1403] = 24'b000000000001001010000100 ; 
		block_ram[1404] = 24'b010000010000000000100000 ; 
		block_ram[1405] = 24'b000000000001001010000010 ; 
		block_ram[1406] = 24'b000000000001001010000001 ; 
		block_ram[1407] = 24'b000000000001001010000000 ; 
		block_ram[1408] = 24'b000000000000010110000000 ; 
		block_ram[1409] = 24'b000000000000010110000001 ; 
		block_ram[1410] = 24'b000000000000010110000010 ; 
		block_ram[1411] = 24'b110000000000000000010000 ; 
		block_ram[1412] = 24'b000000000000010110000100 ; 
		block_ram[1413] = 24'b000000000010100001000000 ; 
		block_ram[1414] = 24'b000000010100000000100000 ; 
		block_ram[1415] = 24'b000000000010100001000010 ; 
		block_ram[1416] = 24'b000000000000010110001000 ; 
		block_ram[1417] = 24'b000000110001000000000000 ; 
		block_ram[1418] = 24'b000100001000000001000000 ; 
		block_ram[1419] = 24'b000000000100111000000000 ; 
		block_ram[1420] = 24'b100010000000001000000000 ; 
		block_ram[1421] = 24'b000000000010100001001000 ; 
		block_ram[1422] = 24'b000000010100000000101000 ; 
		block_ram[1423] = 24'b001001000000000010000000 ; 
		block_ram[1424] = 24'b000000000000010110010000 ; 
		block_ram[1425] = 24'b110000000000000000000010 ; 
		block_ram[1426] = 24'b110000000000000000000001 ; 
		block_ram[1427] = 24'b110000000000000000000000 ; 
		block_ram[1428] = 24'b000101000001000000000000 ; 
		block_ram[1429] = 24'b000000000010100001010000 ; 
		block_ram[1430] = 24'b000000001000101010000000 ; 
		block_ram[1431] = 24'b110000000000000000000100 ; 
		block_ram[1432] = 24'b001000000000100000100000 ; 
		block_ram[1433] = 24'b000000001100000100000100 ; 
		block_ram[1434] = 24'b000000100010010000000100 ; 
		block_ram[1435] = 24'b110000000000000000001000 ; 
		block_ram[1436] = 24'b000000001100000100000001 ; 
		block_ram[1437] = 24'b000000001100000100000000 ; 
		block_ram[1438] = 24'b000000100010010000000000 ; 
		block_ram[1439] = 24'b000000000001001001100000 ; 
		block_ram[1440] = 24'b000000000000010110100000 ; 
		block_ram[1441] = 24'b000001001000001000000000 ; 
		block_ram[1442] = 24'b000000010100000000000100 ; 
		block_ram[1443] = 24'b000000010100000000000101 ; 
		block_ram[1444] = 24'b000000010100000000000010 ; 
		block_ram[1445] = 24'b000000000010100001100000 ; 
		block_ram[1446] = 24'b000000010100000000000000 ; 
		block_ram[1447] = 24'b000000010100000000000001 ; 
		block_ram[1448] = 24'b001000000000100000010000 ; 
		block_ram[1449] = 24'b000000110001000000100000 ; 
		block_ram[1450] = 24'b000000010100000000001100 ; 
		block_ram[1451] = 24'b000010000010000100000000 ; 
		block_ram[1452] = 24'b000000001011000010000000 ; 
		block_ram[1453] = 24'b010100000000010000000000 ; 
		block_ram[1454] = 24'b000000010100000000001000 ; 
		block_ram[1455] = 24'b000000000001001001010000 ; 
		block_ram[1456] = 24'b001000000000100000001000 ; 
		block_ram[1457] = 24'b000000000111010000000000 ; 
		block_ram[1458] = 24'b000000010100000000010100 ; 
		block_ram[1459] = 24'b110000000000000000100000 ; 
		block_ram[1460] = 24'b000000010100000000010010 ; 
		block_ram[1461] = 24'b000010100000000010000000 ; 
		block_ram[1462] = 24'b000000010100000000010000 ; 
		block_ram[1463] = 24'b000000000001001001001000 ; 
		block_ram[1464] = 24'b001000000000100000000000 ; 
		block_ram[1465] = 24'b001000000000100000000001 ; 
		block_ram[1466] = 24'b001000000000100000000010 ; 
		block_ram[1467] = 24'b000000000001001001000100 ; 
		block_ram[1468] = 24'b001000000000100000000100 ; 
		block_ram[1469] = 24'b000000000001001001000010 ; 
		block_ram[1470] = 24'b000000000001001001000001 ; 
		block_ram[1471] = 24'b000000000001001001000000 ; 
		block_ram[1472] = 24'b000000000000010111000000 ; 
		block_ram[1473] = 24'b000000000010100000000100 ; 
		block_ram[1474] = 24'b000100001000000000001000 ; 
		block_ram[1475] = 24'b000000000010100000000110 ; 
		block_ram[1476] = 24'b000000000010100000000001 ; 
		block_ram[1477] = 24'b000000000010100000000000 ; 
		block_ram[1478] = 24'b000000000010100000000011 ; 
		block_ram[1479] = 24'b000000000010100000000010 ; 
		block_ram[1480] = 24'b000100001000000000000010 ; 
		block_ram[1481] = 24'b000000000010100000001100 ; 
		block_ram[1482] = 24'b000100001000000000000000 ; 
		block_ram[1483] = 24'b000100001000000000000001 ; 
		block_ram[1484] = 24'b000000000010100000001001 ; 
		block_ram[1485] = 24'b000000000010100000001000 ; 
		block_ram[1486] = 24'b000100001000000000000100 ; 
		block_ram[1487] = 24'b000000000001001000110000 ; 
		block_ram[1488] = 24'b000000100100001000000000 ; 
		block_ram[1489] = 24'b000000000010100000010100 ; 
		block_ram[1490] = 24'b000000010001110000000000 ; 
		block_ram[1491] = 24'b110000000000000001000000 ; 
		block_ram[1492] = 24'b000000000010100000010001 ; 
		block_ram[1493] = 24'b000000000010100000010000 ; 
		block_ram[1494] = 24'b001010000000000100000000 ; 
		block_ram[1495] = 24'b000000000001001000101000 ; 
		block_ram[1496] = 24'b000000100100001000001000 ; 
		block_ram[1497] = 24'b000011000000010000000000 ; 
		block_ram[1498] = 24'b000100001000000000010000 ; 
		block_ram[1499] = 24'b000000000001001000100100 ; 
		block_ram[1500] = 24'b010000010000000010000000 ; 
		block_ram[1501] = 24'b000000000001001000100010 ; 
		block_ram[1502] = 24'b000000000001001000100001 ; 
		block_ram[1503] = 24'b000000000001001000100000 ; 
		block_ram[1504] = 24'b010010000001000000000000 ; 
		block_ram[1505] = 24'b000000000010100000100100 ; 
		block_ram[1506] = 24'b000000010100000001000100 ; 
		block_ram[1507] = 24'b001000100000010000000000 ; 
		block_ram[1508] = 24'b000000000010100000100001 ; 
		block_ram[1509] = 24'b000000000010100000100000 ; 
		block_ram[1510] = 24'b000000010100000001000000 ; 
		block_ram[1511] = 24'b000000000001001000011000 ; 
		block_ram[1512] = 24'b000000010010011000000000 ; 
		block_ram[1513] = 24'b100000000100000010000000 ; 
		block_ram[1514] = 24'b000100001000000000100000 ; 
		block_ram[1515] = 24'b000000000001001000010100 ; 
		block_ram[1516] = 24'b000001100000000100000000 ; 
		block_ram[1517] = 24'b000000000001001000010010 ; 
		block_ram[1518] = 24'b000000000001001000010001 ; 
		block_ram[1519] = 24'b000000000001001000010000 ; 
		block_ram[1520] = 24'b000000100100001000100000 ; 
		block_ram[1521] = 24'b000100010000000100000000 ; 
		block_ram[1522] = 24'b000001000010000010000000 ; 
		block_ram[1523] = 24'b000000000001001000001100 ; 
		block_ram[1524] = 24'b100000001000010000000000 ; 
		block_ram[1525] = 24'b000000000001001000001010 ; 
		block_ram[1526] = 24'b000000000001001000001001 ; 
		block_ram[1527] = 24'b000000000001001000001000 ; 
		block_ram[1528] = 24'b001000000000100001000000 ; 
		block_ram[1529] = 24'b000000000001001000000110 ; 
		block_ram[1530] = 24'b000000000001001000000101 ; 
		block_ram[1531] = 24'b000000000001001000000100 ; 
		block_ram[1532] = 24'b000000000001001000000011 ; 
		block_ram[1533] = 24'b000000000001001000000010 ; 
		block_ram[1534] = 24'b000000000001001000000001 ; 
		block_ram[1535] = 24'b000000000001001000000000 ; 
		block_ram[1536] = 24'b000000000000011000000000 ; 
		block_ram[1537] = 24'b000000000000011000000001 ; 
		block_ram[1538] = 24'b000000000000011000000010 ; 
		block_ram[1539] = 24'b000000000000011000000011 ; 
		block_ram[1540] = 24'b000000000000011000000100 ; 
		block_ram[1541] = 24'b000000000000011000000101 ; 
		block_ram[1542] = 24'b000000000000011000000110 ; 
		block_ram[1543] = 24'b000100100000000010000000 ; 
		block_ram[1544] = 24'b000000000000011000001000 ; 
		block_ram[1545] = 24'b000000000000011000001001 ; 
		block_ram[1546] = 24'b000000000000011000001010 ; 
		block_ram[1547] = 24'b100000001001000000000000 ; 
		block_ram[1548] = 24'b000000000000011000001100 ; 
		block_ram[1549] = 24'b000000010000100000100000 ; 
		block_ram[1550] = 24'b000000000110000001000000 ; 
		block_ram[1551] = 24'b000000000110000001000001 ; 
		block_ram[1552] = 24'b000000000000011000010000 ; 
		block_ram[1553] = 24'b000000000000011000010001 ; 
		block_ram[1554] = 24'b000000000000011000010010 ; 
		block_ram[1555] = 24'b001000000100000000100000 ; 
		block_ram[1556] = 24'b000000000000011000010100 ; 
		block_ram[1557] = 24'b100001000000000001000000 ; 
		block_ram[1558] = 24'b000000001000100100000000 ; 
		block_ram[1559] = 24'b000000001000100100000001 ; 
		block_ram[1560] = 24'b000000000000011000011000 ; 
		block_ram[1561] = 24'b000100000010000100000000 ; 
		block_ram[1562] = 24'b000001010000000010000000 ; 
		block_ram[1563] = 24'b000000100000101001000000 ; 
		block_ram[1564] = 24'b001000100001000000000000 ; 
		block_ram[1565] = 24'b000000001100001010000000 ; 
		block_ram[1566] = 24'b000000000110000001010000 ; 
		block_ram[1567] = 24'b010010000000010000000000 ; 
		block_ram[1568] = 24'b000000000000011000100000 ; 
		block_ram[1569] = 24'b000000000000011000100001 ; 
		block_ram[1570] = 24'b000000000000011000100010 ; 
		block_ram[1571] = 24'b001000000100000000010000 ; 
		block_ram[1572] = 24'b000000000000011000100100 ; 
		block_ram[1573] = 24'b000000010000100000001000 ; 
		block_ram[1574] = 24'b000011000001000000000000 ; 
		block_ram[1575] = 24'b000000010000100000001010 ; 
		block_ram[1576] = 24'b000000000000011000101000 ; 
		block_ram[1577] = 24'b000000010000100000000100 ; 
		block_ram[1578] = 24'b010000100000000100000000 ; 
		block_ram[1579] = 24'b000000010000100000000110 ; 
		block_ram[1580] = 24'b000000010000100000000001 ; 
		block_ram[1581] = 24'b000000010000100000000000 ; 
		block_ram[1582] = 24'b000000000110000001100000 ; 
		block_ram[1583] = 24'b000000010000100000000010 ; 
		block_ram[1584] = 24'b000000000000011000110000 ; 
		block_ram[1585] = 24'b001000000100000000000010 ; 
		block_ram[1586] = 24'b001000000100000000000001 ; 
		block_ram[1587] = 24'b001000000100000000000000 ; 
		block_ram[1588] = 24'b010000000010000010000000 ; 
		block_ram[1589] = 24'b000000010000100000011000 ; 
		block_ram[1590] = 24'b000000001000100100100000 ; 
		block_ram[1591] = 24'b001000000100000000000100 ; 
		block_ram[1592] = 24'b000010001000000001000000 ; 
		block_ram[1593] = 24'b000000010000100000010100 ; 
		block_ram[1594] = 24'b000000000011110000000000 ; 
		block_ram[1595] = 24'b001000000100000000001000 ; 
		block_ram[1596] = 24'b000000010000100000010001 ; 
		block_ram[1597] = 24'b000000010000100000010000 ; 
		block_ram[1598] = 24'b100100000000001000000000 ; 
		block_ram[1599] = 24'b000000000001000111000000 ; 
		block_ram[1600] = 24'b000000000000011001000000 ; 
		block_ram[1601] = 24'b000000000000011001000001 ; 
		block_ram[1602] = 24'b000000000000011001000010 ; 
		block_ram[1603] = 24'b000010010000000100000000 ; 
		block_ram[1604] = 24'b000000000000011001000100 ; 
		block_ram[1605] = 24'b100001000000000000010000 ; 
		block_ram[1606] = 24'b000000000110000000001000 ; 
		block_ram[1607] = 24'b000000000110000000001001 ; 
		block_ram[1608] = 24'b000000000000011001001000 ; 
		block_ram[1609] = 24'b011000000000000010000000 ; 
		block_ram[1610] = 24'b000000000110000000000100 ; 
		block_ram[1611] = 24'b000000000110000000000101 ; 
		block_ram[1612] = 24'b000000000110000000000010 ; 
		block_ram[1613] = 24'b000000000110000000000011 ; 
		block_ram[1614] = 24'b000000000110000000000000 ; 
		block_ram[1615] = 24'b000000000110000000000001 ; 
		block_ram[1616] = 24'b000000000000011001010000 ; 
		block_ram[1617] = 24'b100001000000000000000100 ; 
		block_ram[1618] = 24'b010100000001000000000000 ; 
		block_ram[1619] = 24'b000000001010010010000000 ; 
		block_ram[1620] = 24'b100001000000000000000001 ; 
		block_ram[1621] = 24'b100001000000000000000000 ; 
		block_ram[1622] = 24'b000000000110000000011000 ; 
		block_ram[1623] = 24'b100001000000000000000010 ; 
		block_ram[1624] = 24'b000010001000000000100000 ; 
		block_ram[1625] = 24'b000000010101010000000000 ; 
		block_ram[1626] = 24'b000000000110000000010100 ; 
		block_ram[1627] = 24'b000000100000101000000000 ; 
		block_ram[1628] = 24'b000000000110000000010010 ; 
		block_ram[1629] = 24'b100001000000000000001000 ; 
		block_ram[1630] = 24'b000000000110000000010000 ; 
		block_ram[1631] = 24'b000000000001000110100000 ; 
		block_ram[1632] = 24'b000000000000011001100000 ; 
		block_ram[1633] = 24'b000000100011000000000000 ; 
		block_ram[1634] = 24'b100000000000100010000000 ; 
		block_ram[1635] = 24'b000000100011000000000010 ; 
		block_ram[1636] = 24'b001100000000000100000000 ; 
		block_ram[1637] = 24'b000000010000100001001000 ; 
		block_ram[1638] = 24'b000000000110000000101000 ; 
		block_ram[1639] = 24'b010000001000001000000000 ; 
		block_ram[1640] = 24'b000010001000000000010000 ; 
		block_ram[1641] = 24'b000000010000100001000100 ; 
		block_ram[1642] = 24'b000000000110000000100100 ; 
		block_ram[1643] = 24'b000101000000010000000000 ; 
		block_ram[1644] = 24'b000000000110000000100010 ; 
		block_ram[1645] = 24'b000000010000100001000000 ; 
		block_ram[1646] = 24'b000000000110000000100000 ; 
		block_ram[1647] = 24'b000000000001000110010000 ; 
		block_ram[1648] = 24'b000010001000000000001000 ; 
		block_ram[1649] = 24'b000000100011000000010000 ; 
		block_ram[1650] = 24'b000000110000010000000100 ; 
		block_ram[1651] = 24'b001000000100000001000000 ; 
		block_ram[1652] = 24'b000000000101101000000000 ; 
		block_ram[1653] = 24'b100001000000000000100000 ; 
		block_ram[1654] = 24'b000000110000010000000000 ; 
		block_ram[1655] = 24'b000000000001000110001000 ; 
		block_ram[1656] = 24'b000010001000000000000000 ; 
		block_ram[1657] = 24'b000010001000000000000001 ; 
		block_ram[1658] = 24'b000010001000000000000010 ; 
		block_ram[1659] = 24'b000000000001000110000100 ; 
		block_ram[1660] = 24'b000010001000000000000100 ; 
		block_ram[1661] = 24'b000000000001000110000010 ; 
		block_ram[1662] = 24'b000000000001000110000001 ; 
		block_ram[1663] = 24'b000000000001000110000000 ; 
		block_ram[1664] = 24'b000000000000011010000000 ; 
		block_ram[1665] = 24'b000000000000011010000001 ; 
		block_ram[1666] = 24'b000000000000011010000010 ; 
		block_ram[1667] = 24'b000100100000000000000100 ; 
		block_ram[1668] = 24'b000000000000011010000100 ; 
		block_ram[1669] = 24'b000100100000000000000010 ; 
		block_ram[1670] = 24'b000100100000000000000001 ; 
		block_ram[1671] = 24'b000100100000000000000000 ; 
		block_ram[1672] = 24'b000000000000011010001000 ; 
		block_ram[1673] = 24'b011000000000000001000000 ; 
		block_ram[1674] = 24'b000001010000000000010000 ; 
		block_ram[1675] = 24'b000000000100110100000000 ; 
		block_ram[1676] = 24'b100010000000000100000000 ; 
		block_ram[1677] = 24'b000000001100001000010000 ; 
		block_ram[1678] = 24'b000000000110000011000000 ; 
		block_ram[1679] = 24'b000100100000000000001000 ; 
		block_ram[1680] = 24'b000000000000011010010000 ; 
		block_ram[1681] = 24'b000010000001100000000000 ; 
		block_ram[1682] = 24'b000001010000000000001000 ; 
		block_ram[1683] = 24'b000000001010010001000000 ; 
		block_ram[1684] = 24'b010000000010000000100000 ; 
		block_ram[1685] = 24'b000000001100001000001000 ; 
		block_ram[1686] = 24'b000000001000100110000000 ; 
		block_ram[1687] = 24'b000100100000000000010000 ; 
		block_ram[1688] = 24'b000001010000000000000010 ; 
		block_ram[1689] = 24'b000000001100001000000100 ; 
		block_ram[1690] = 24'b000001010000000000000000 ; 
		block_ram[1691] = 24'b000001010000000000000001 ; 
		block_ram[1692] = 24'b000000001100001000000001 ; 
		block_ram[1693] = 24'b000000001100001000000000 ; 
		block_ram[1694] = 24'b000001010000000000000100 ; 
		block_ram[1695] = 24'b000000000001000101100000 ; 
		block_ram[1696] = 24'b000000000000011010100000 ; 
		block_ram[1697] = 24'b000001001000000100000000 ; 
		block_ram[1698] = 24'b100000000000100001000000 ; 
		block_ram[1699] = 24'b000001001000000100000010 ; 
		block_ram[1700] = 24'b010000000010000000010000 ; 
		block_ram[1701] = 24'b000000010000100010001000 ; 
		block_ram[1702] = 24'b000000010100001100000000 ; 
		block_ram[1703] = 24'b000100100000000000100000 ; 
		block_ram[1704] = 24'b000100000101000000000000 ; 
		block_ram[1705] = 24'b000000010000100010000100 ; 
		block_ram[1706] = 24'b000001010000000000110000 ; 
		block_ram[1707] = 24'b000010000010001000000000 ; 
		block_ram[1708] = 24'b000000010000100010000001 ; 
		block_ram[1709] = 24'b000000010000100010000000 ; 
		block_ram[1710] = 24'b001000001000010000000000 ; 
		block_ram[1711] = 24'b000000000001000101010000 ; 
		block_ram[1712] = 24'b010000000010000000000100 ; 
		block_ram[1713] = 24'b000001001000000100010000 ; 
		block_ram[1714] = 24'b000000101001001000000000 ; 
		block_ram[1715] = 24'b001000000100000010000000 ; 
		block_ram[1716] = 24'b010000000010000000000000 ; 
		block_ram[1717] = 24'b010000000010000000000001 ; 
		block_ram[1718] = 24'b010000000010000000000010 ; 
		block_ram[1719] = 24'b000000000001000101001000 ; 
		block_ram[1720] = 24'b000001010000000000100010 ; 
		block_ram[1721] = 24'b100000100000010000000000 ; 
		block_ram[1722] = 24'b000001010000000000100000 ; 
		block_ram[1723] = 24'b000000000001000101000100 ; 
		block_ram[1724] = 24'b010000000010000000001000 ; 
		block_ram[1725] = 24'b000000000001000101000010 ; 
		block_ram[1726] = 24'b000000000001000101000001 ; 
		block_ram[1727] = 24'b000000000001000101000000 ; 
		block_ram[1728] = 24'b000000000000011011000000 ; 
		block_ram[1729] = 24'b011000000000000000001000 ; 
		block_ram[1730] = 24'b100000000000100000100000 ; 
		block_ram[1731] = 24'b000000001010010000010000 ; 
		block_ram[1732] = 24'b000000011001000000000000 ; 
		block_ram[1733] = 24'b000000000010101100000000 ; 
		block_ram[1734] = 24'b000000000110000010001000 ; 
		block_ram[1735] = 24'b000100100000000001000000 ; 
		block_ram[1736] = 24'b011000000000000000000001 ; 
		block_ram[1737] = 24'b011000000000000000000000 ; 
		block_ram[1738] = 24'b000000000110000010000100 ; 
		block_ram[1739] = 24'b011000000000000000000010 ; 
		block_ram[1740] = 24'b000000000110000010000010 ; 
		block_ram[1741] = 24'b011000000000000000000100 ; 
		block_ram[1742] = 24'b000000000110000010000000 ; 
		block_ram[1743] = 24'b000000000001000100110000 ; 
		block_ram[1744] = 24'b000000100100000100000000 ; 
		block_ram[1745] = 24'b000000001010010000000010 ; 
		block_ram[1746] = 24'b000000001010010000000001 ; 
		block_ram[1747] = 24'b000000001010010000000000 ; 
		block_ram[1748] = 24'b000000011001000000010000 ; 
		block_ram[1749] = 24'b100001000000000010000000 ; 
		block_ram[1750] = 24'b001010000000001000000000 ; 
		block_ram[1751] = 24'b000000000001000100101000 ; 
		block_ram[1752] = 24'b000000100100000100001000 ; 
		block_ram[1753] = 24'b011000000000000000010000 ; 
		block_ram[1754] = 24'b000001010000000001000000 ; 
		block_ram[1755] = 24'b000000000001000100100100 ; 
		block_ram[1756] = 24'b000100000000110000000000 ; 
		block_ram[1757] = 24'b000000000001000100100010 ; 
		block_ram[1758] = 24'b000000000001000100100001 ; 
		block_ram[1759] = 24'b000000000001000100100000 ; 
		block_ram[1760] = 24'b100000000000100000000010 ; 
		block_ram[1761] = 24'b000000100011000010000000 ; 
		block_ram[1762] = 24'b100000000000100000000000 ; 
		block_ram[1763] = 24'b100000000000100000000001 ; 
		block_ram[1764] = 24'b000000011001000000100000 ; 
		block_ram[1765] = 24'b000010000100010000000000 ; 
		block_ram[1766] = 24'b100000000000100000000100 ; 
		block_ram[1767] = 24'b000000000001000100011000 ; 
		block_ram[1768] = 24'b000000010010010100000000 ; 
		block_ram[1769] = 24'b011000000000000000100000 ; 
		block_ram[1770] = 24'b100000000000100000001000 ; 
		block_ram[1771] = 24'b000000000001000100010100 ; 
		block_ram[1772] = 24'b000001100000001000000000 ; 
		block_ram[1773] = 24'b000000000001000100010010 ; 
		block_ram[1774] = 24'b000000000001000100010001 ; 
		block_ram[1775] = 24'b000000000001000100010000 ; 
		block_ram[1776] = 24'b000000100100000100100000 ; 
		block_ram[1777] = 24'b000100010000001000000000 ; 
		block_ram[1778] = 24'b100000000000100000010000 ; 
		block_ram[1779] = 24'b000000000001000100001100 ; 
		block_ram[1780] = 24'b010000000010000001000000 ; 
		block_ram[1781] = 24'b000000000001000100001010 ; 
		block_ram[1782] = 24'b000000000001000100001001 ; 
		block_ram[1783] = 24'b000000000001000100001000 ; 
		block_ram[1784] = 24'b000010001000000010000000 ; 
		block_ram[1785] = 24'b000000000001000100000110 ; 
		block_ram[1786] = 24'b000000000001000100000101 ; 
		block_ram[1787] = 24'b000000000001000100000100 ; 
		block_ram[1788] = 24'b000000000001000100000011 ; 
		block_ram[1789] = 24'b000000000001000100000010 ; 
		block_ram[1790] = 24'b000000000001000100000001 ; 
		block_ram[1791] = 24'b000000000001000100000000 ; 
		block_ram[1792] = 24'b000000000000011100000000 ; 
		block_ram[1793] = 24'b000000000000011100000001 ; 
		block_ram[1794] = 24'b000000000000011100000010 ; 
		block_ram[1795] = 24'b000010010000000001000000 ; 
		block_ram[1796] = 24'b000000000000011100000100 ; 
		block_ram[1797] = 24'b010000000101000000000000 ; 
		block_ram[1798] = 24'b000000001000100000010000 ; 
		block_ram[1799] = 24'b000000001000100000010001 ; 
		block_ram[1800] = 24'b000000000000011100001000 ; 
		block_ram[1801] = 24'b000100000010000000010000 ; 
		block_ram[1802] = 24'b010000100000000000100000 ; 
		block_ram[1803] = 24'b000000000100110010000000 ; 
		block_ram[1804] = 24'b100010000000000010000000 ; 
		block_ram[1805] = 24'b000000010000100100100000 ; 
		block_ram[1806] = 24'b000000000110000101000000 ; 
		block_ram[1807] = 24'b001001000000001000000000 ; 
		block_ram[1808] = 24'b000000000000011100010000 ; 
		block_ram[1809] = 24'b000100000010000000001000 ; 
		block_ram[1810] = 24'b000000001000100000000100 ; 
		block_ram[1811] = 24'b000000001000100000000101 ; 
		block_ram[1812] = 24'b000000001000100000000010 ; 
		block_ram[1813] = 24'b000000001000100000000011 ; 
		block_ram[1814] = 24'b000000001000100000000000 ; 
		block_ram[1815] = 24'b000000001000100000000001 ; 
		block_ram[1816] = 24'b000100000010000000000001 ; 
		block_ram[1817] = 24'b000100000010000000000000 ; 
		block_ram[1818] = 24'b000000001000100000001100 ; 
		block_ram[1819] = 24'b000100000010000000000010 ; 
		block_ram[1820] = 24'b000000001000100000001010 ; 
		block_ram[1821] = 24'b000100000010000000000100 ; 
		block_ram[1822] = 24'b000000001000100000001000 ; 
		block_ram[1823] = 24'b000000000001000011100000 ; 
		block_ram[1824] = 24'b000000000000011100100000 ; 
		block_ram[1825] = 24'b000001001000000010000000 ; 
		block_ram[1826] = 24'b010000100000000000001000 ; 
		block_ram[1827] = 24'b000001001000000010000010 ; 
		block_ram[1828] = 24'b001100000000000001000000 ; 
		block_ram[1829] = 24'b000000010000100100001000 ; 
		block_ram[1830] = 24'b000000001000100000110000 ; 
		block_ram[1831] = 24'b100000000010010000000000 ; 
		block_ram[1832] = 24'b010000100000000000000010 ; 
		block_ram[1833] = 24'b000000010000100100000100 ; 
		block_ram[1834] = 24'b010000100000000000000000 ; 
		block_ram[1835] = 24'b010000100000000000000001 ; 
		block_ram[1836] = 24'b000000001011001000000000 ; 
		block_ram[1837] = 24'b000000010000100100000000 ; 
		block_ram[1838] = 24'b010000100000000000000100 ; 
		block_ram[1839] = 24'b000000000001000011010000 ; 
		block_ram[1840] = 24'b100000010001000000000000 ; 
		block_ram[1841] = 24'b000001001000000010010000 ; 
		block_ram[1842] = 24'b000000001000100000100100 ; 
		block_ram[1843] = 24'b001000000100000100000000 ; 
		block_ram[1844] = 24'b000000001000100000100010 ; 
		block_ram[1845] = 24'b000010100000001000000000 ; 
		block_ram[1846] = 24'b000000001000100000100000 ; 
		block_ram[1847] = 24'b000000000001000011001000 ; 
		block_ram[1848] = 24'b000001000100010000000100 ; 
		block_ram[1849] = 24'b000100000010000000100000 ; 
		block_ram[1850] = 24'b010000100000000000010000 ; 
		block_ram[1851] = 24'b000000000001000011000100 ; 
		block_ram[1852] = 24'b000001000100010000000000 ; 
		block_ram[1853] = 24'b000000000001000011000010 ; 
		block_ram[1854] = 24'b000000000001000011000001 ; 
		block_ram[1855] = 24'b000000000001000011000000 ; 
		block_ram[1856] = 24'b000000000000011101000000 ; 
		block_ram[1857] = 24'b000010010000000000000010 ; 
		block_ram[1858] = 24'b000010010000000000000001 ; 
		block_ram[1859] = 24'b000010010000000000000000 ; 
		block_ram[1860] = 24'b001100000000000000100000 ; 
		block_ram[1861] = 24'b000000000010101010000000 ; 
		block_ram[1862] = 24'b000000000110000100001000 ; 
		block_ram[1863] = 24'b000010010000000000000100 ; 
		block_ram[1864] = 24'b000001000001100000000000 ; 
		block_ram[1865] = 24'b000000101000010000000100 ; 
		block_ram[1866] = 24'b000000000110000100000100 ; 
		block_ram[1867] = 24'b000010010000000000001000 ; 
		block_ram[1868] = 24'b000000000110000100000010 ; 
		block_ram[1869] = 24'b000000101000010000000000 ; 
		block_ram[1870] = 24'b000000000110000100000000 ; 
		block_ram[1871] = 24'b000000000001000010110000 ; 
		block_ram[1872] = 24'b000000100100000010000000 ; 
		block_ram[1873] = 24'b000000100100000010000001 ; 
		block_ram[1874] = 24'b000000001000100001000100 ; 
		block_ram[1875] = 24'b000010010000000000010000 ; 
		block_ram[1876] = 24'b000000001000100001000010 ; 
		block_ram[1877] = 24'b100001000000000100000000 ; 
		block_ram[1878] = 24'b000000001000100001000000 ; 
		block_ram[1879] = 24'b000000000001000010101000 ; 
		block_ram[1880] = 24'b000000100100000010001000 ; 
		block_ram[1881] = 24'b000100000010000001000000 ; 
		block_ram[1882] = 24'b101000000000010000000000 ; 
		block_ram[1883] = 24'b000000000001000010100100 ; 
		block_ram[1884] = 24'b010000010000001000000000 ; 
		block_ram[1885] = 24'b000000000001000010100010 ; 
		block_ram[1886] = 24'b000000000001000010100001 ; 
		block_ram[1887] = 24'b000000000001000010100000 ; 
		block_ram[1888] = 24'b001100000000000000000100 ; 
		block_ram[1889] = 24'b000000100011000100000000 ; 
		block_ram[1890] = 24'b000000001101010000000000 ; 
		block_ram[1891] = 24'b000010010000000000100000 ; 
		block_ram[1892] = 24'b001100000000000000000000 ; 
		block_ram[1893] = 24'b001100000000000000000001 ; 
		block_ram[1894] = 24'b001100000000000000000010 ; 
		block_ram[1895] = 24'b000000000001000010011000 ; 
		block_ram[1896] = 24'b000000010010010010000000 ; 
		block_ram[1897] = 24'b100000000100001000000000 ; 
		block_ram[1898] = 24'b010000100000000001000000 ; 
		block_ram[1899] = 24'b000000000001000010010100 ; 
		block_ram[1900] = 24'b001100000000000000001000 ; 
		block_ram[1901] = 24'b000000000001000010010010 ; 
		block_ram[1902] = 24'b000000000001000010010001 ; 
		block_ram[1903] = 24'b000000000001000010010000 ; 
		block_ram[1904] = 24'b000000100100000010100000 ; 
		block_ram[1905] = 24'b010000000000110000000000 ; 
		block_ram[1906] = 24'b000001000010001000000000 ; 
		block_ram[1907] = 24'b000000000001000010001100 ; 
		block_ram[1908] = 24'b001100000000000000010000 ; 
		block_ram[1909] = 24'b000000000001000010001010 ; 
		block_ram[1910] = 24'b000000000001000010001001 ; 
		block_ram[1911] = 24'b000000000001000010001000 ; 
		block_ram[1912] = 24'b000010001000000100000000 ; 
		block_ram[1913] = 24'b000000000001000010000110 ; 
		block_ram[1914] = 24'b000000000001000010000101 ; 
		block_ram[1915] = 24'b000000000001000010000100 ; 
		block_ram[1916] = 24'b000000000001000010000011 ; 
		block_ram[1917] = 24'b000000000001000010000010 ; 
		block_ram[1918] = 24'b000000000001000010000001 ; 
		block_ram[1919] = 24'b000000000001000010000000 ; 
		block_ram[1920] = 24'b000000000000011110000000 ; 
		block_ram[1921] = 24'b000001001000000000100000 ; 
		block_ram[1922] = 24'b001000000011000000000000 ; 
		block_ram[1923] = 24'b000000000100110000001000 ; 
		block_ram[1924] = 24'b100010000000000000001000 ; 
		block_ram[1925] = 24'b000000000010101001000000 ; 
		block_ram[1926] = 24'b000000001000100010010000 ; 
		block_ram[1927] = 24'b000100100000000100000000 ; 
		block_ram[1928] = 24'b100010000000000000000100 ; 
		block_ram[1929] = 24'b000000000100110000000010 ; 
		block_ram[1930] = 24'b000000000100110000000001 ; 
		block_ram[1931] = 24'b000000000100110000000000 ; 
		block_ram[1932] = 24'b100010000000000000000000 ; 
		block_ram[1933] = 24'b100010000000000000000001 ; 
		block_ram[1934] = 24'b100010000000000000000010 ; 
		block_ram[1935] = 24'b000000000001000001110000 ; 
		block_ram[1936] = 24'b000000100100000001000000 ; 
		block_ram[1937] = 24'b000000100100000001000001 ; 
		block_ram[1938] = 24'b000000001000100010000100 ; 
		block_ram[1939] = 24'b110000000000001000000000 ; 
		block_ram[1940] = 24'b000000001000100010000010 ; 
		block_ram[1941] = 24'b001000010000010000000000 ; 
		block_ram[1942] = 24'b000000001000100010000000 ; 
		block_ram[1943] = 24'b000000000001000001101000 ; 
		block_ram[1944] = 24'b000000100100000001001000 ; 
		block_ram[1945] = 24'b000100000010000010000000 ; 
		block_ram[1946] = 24'b000001010000000100000000 ; 
		block_ram[1947] = 24'b000000000001000001100100 ; 
		block_ram[1948] = 24'b100010000000000000010000 ; 
		block_ram[1949] = 24'b000000000001000001100010 ; 
		block_ram[1950] = 24'b000000000001000001100001 ; 
		block_ram[1951] = 24'b000000000001000001100000 ; 
		block_ram[1952] = 24'b000001001000000000000001 ; 
		block_ram[1953] = 24'b000001001000000000000000 ; 
		block_ram[1954] = 24'b000000010100001000000100 ; 
		block_ram[1955] = 24'b000001001000000000000010 ; 
		block_ram[1956] = 24'b000000010100001000000010 ; 
		block_ram[1957] = 24'b000001001000000000000100 ; 
		block_ram[1958] = 24'b000000010100001000000000 ; 
		block_ram[1959] = 24'b000000000001000001011000 ; 
		block_ram[1960] = 24'b000000010010010001000000 ; 
		block_ram[1961] = 24'b000001001000000000001000 ; 
		block_ram[1962] = 24'b010000100000000010000000 ; 
		block_ram[1963] = 24'b000000000001000001010100 ; 
		block_ram[1964] = 24'b100010000000000000100000 ; 
		block_ram[1965] = 24'b000000000001000001010010 ; 
		block_ram[1966] = 24'b000000000001000001010001 ; 
		block_ram[1967] = 24'b000000000001000001010000 ; 
		block_ram[1968] = 24'b000000100100000001100000 ; 
		block_ram[1969] = 24'b000001001000000000010000 ; 
		block_ram[1970] = 24'b000110000000010000000000 ; 
		block_ram[1971] = 24'b000000000001000001001100 ; 
		block_ram[1972] = 24'b010000000010000100000000 ; 
		block_ram[1973] = 24'b000000000001000001001010 ; 
		block_ram[1974] = 24'b000000000001000001001001 ; 
		block_ram[1975] = 24'b000000000001000001001000 ; 
		block_ram[1976] = 24'b001000000000101000000000 ; 
		block_ram[1977] = 24'b000000000001000001000110 ; 
		block_ram[1978] = 24'b000000000001000001000101 ; 
		block_ram[1979] = 24'b000000000001000001000100 ; 
		block_ram[1980] = 24'b000000000001000001000011 ; 
		block_ram[1981] = 24'b000000000001000001000010 ; 
		block_ram[1982] = 24'b000000000001000001000001 ; 
		block_ram[1983] = 24'b000000000001000001000000 ; 
		block_ram[1984] = 24'b000000100100000000010000 ; 
		block_ram[1985] = 24'b000000000010101000000100 ; 
		block_ram[1986] = 24'b000000100100000000010010 ; 
		block_ram[1987] = 24'b000010010000000010000000 ; 
		block_ram[1988] = 24'b000000000010101000000001 ; 
		block_ram[1989] = 24'b000000000010101000000000 ; 
		block_ram[1990] = 24'b010001000000010000000000 ; 
		block_ram[1991] = 24'b000000000001000000111000 ; 
		block_ram[1992] = 24'b000000010010010000100000 ; 
		block_ram[1993] = 24'b011000000000000100000000 ; 
		block_ram[1994] = 24'b000100001000001000000000 ; 
		block_ram[1995] = 24'b000000000001000000110100 ; 
		block_ram[1996] = 24'b100010000000000001000000 ; 
		block_ram[1997] = 24'b000000000001000000110010 ; 
		block_ram[1998] = 24'b000000000001000000110001 ; 
		block_ram[1999] = 24'b000000000001000000110000 ; 
		block_ram[2000] = 24'b000000100100000000000000 ; 
		block_ram[2001] = 24'b000000100100000000000001 ; 
		block_ram[2002] = 24'b000000100100000000000010 ; 
		block_ram[2003] = 24'b000000000001000000101100 ; 
		block_ram[2004] = 24'b000000100100000000000100 ; 
		block_ram[2005] = 24'b000000000001000000101010 ; 
		block_ram[2006] = 24'b000000000001000000101001 ; 
		block_ram[2007] = 24'b000000000001000000101000 ; 
		block_ram[2008] = 24'b000000100100000000001000 ; 
		block_ram[2009] = 24'b000000000001000000100110 ; 
		block_ram[2010] = 24'b000000000001000000100101 ; 
		block_ram[2011] = 24'b000000000001000000100100 ; 
		block_ram[2012] = 24'b000000000001000000100011 ; 
		block_ram[2013] = 24'b000000000001000000100010 ; 
		block_ram[2014] = 24'b000000000001000000100001 ; 
		block_ram[2015] = 24'b000000000001000000100000 ; 
		block_ram[2016] = 24'b000000010010010000001000 ; 
		block_ram[2017] = 24'b000001001000000001000000 ; 
		block_ram[2018] = 24'b100000000000100100000000 ; 
		block_ram[2019] = 24'b000000000001000000011100 ; 
		block_ram[2020] = 24'b001100000000000010000000 ; 
		block_ram[2021] = 24'b000000000001000000011010 ; 
		block_ram[2022] = 24'b000000000001000000011001 ; 
		block_ram[2023] = 24'b000000000001000000011000 ; 
		block_ram[2024] = 24'b000000010010010000000000 ; 
		block_ram[2025] = 24'b000000000001000000010110 ; 
		block_ram[2026] = 24'b000000000001000000010101 ; 
		block_ram[2027] = 24'b000000000001000000010100 ; 
		block_ram[2028] = 24'b000000000001000000010011 ; 
		block_ram[2029] = 24'b000000000001000000010010 ; 
		block_ram[2030] = 24'b000000000001000000010001 ; 
		block_ram[2031] = 24'b000000000001000000010000 ; 
		block_ram[2032] = 24'b000000100100000000100000 ; 
		block_ram[2033] = 24'b000000000001000000001110 ; 
		block_ram[2034] = 24'b000000000001000000001101 ; 
		block_ram[2035] = 24'b000000000001000000001100 ; 
		block_ram[2036] = 24'b000000000001000000001011 ; 
		block_ram[2037] = 24'b000000000001000000001010 ; 
		block_ram[2038] = 24'b000000000001000000001001 ; 
		block_ram[2039] = 24'b000000000001000000001000 ; 
		block_ram[2040] = 24'b000000000001000000000111 ; 
		block_ram[2041] = 24'b000000000001000000000110 ; 
		block_ram[2042] = 24'b000000000001000000000101 ; 
		block_ram[2043] = 24'b000000000001000000000100 ; 
		block_ram[2044] = 24'b000000000001000000000011 ; 
		block_ram[2045] = 24'b000000000001000000000010 ; 
		block_ram[2046] = 24'b000000000001000000000001 ; 
		block_ram[2047] = 24'b000000000001000000000000 ; 
		block_ram[2048] = 24'b000000000000100000000000 ; 
		block_ram[2049] = 24'b000000000000100000000001 ; 
		block_ram[2050] = 24'b000000000000100000000010 ; 
		block_ram[2051] = 24'b000000000000100000000011 ; 
		block_ram[2052] = 24'b000000000000100000000100 ; 
		block_ram[2053] = 24'b000000000000100000000101 ; 
		block_ram[2054] = 24'b000000000000100000000110 ; 
		block_ram[2055] = 24'b000000000000100000000111 ; 
		block_ram[2056] = 24'b000000000000100000001000 ; 
		block_ram[2057] = 24'b000000000000100000001001 ; 
		block_ram[2058] = 24'b000000000000100000001010 ; 
		block_ram[2059] = 24'b000000000000100000001011 ; 
		block_ram[2060] = 24'b000000000000100000001100 ; 
		block_ram[2061] = 24'b000000000000100000001101 ; 
		block_ram[2062] = 24'b000000000000100000001110 ; 
		block_ram[2063] = 24'b000100001010000000000000 ; 
		block_ram[2064] = 24'b000000000000100000010000 ; 
		block_ram[2065] = 24'b000000000000100000010001 ; 
		block_ram[2066] = 24'b000000000000100000010010 ; 
		block_ram[2067] = 24'b000000000000100000010011 ; 
		block_ram[2068] = 24'b000000000000100000010100 ; 
		block_ram[2069] = 24'b000000000000100000010101 ; 
		block_ram[2070] = 24'b000000000000100000010110 ; 
		block_ram[2071] = 24'b000001000000000010100000 ; 
		block_ram[2072] = 24'b000000000000100000011000 ; 
		block_ram[2073] = 24'b000000000000100000011001 ; 
		block_ram[2074] = 24'b000000000000100000011010 ; 
		block_ram[2075] = 24'b000000100000010001000000 ; 
		block_ram[2076] = 24'b000000000000100000011100 ; 
		block_ram[2077] = 24'b100000000001000100000000 ; 
		block_ram[2078] = 24'b001000010100000000000000 ; 
		block_ram[2079] = 24'b000000100000010001000100 ; 
		block_ram[2080] = 24'b000000000000100000100000 ; 
		block_ram[2081] = 24'b000000000000100000100001 ; 
		block_ram[2082] = 24'b000000000000100000100010 ; 
		block_ram[2083] = 24'b000000000000100000100011 ; 
		block_ram[2084] = 24'b000000000000100000100100 ; 
		block_ram[2085] = 24'b000000000000100000100101 ; 
		block_ram[2086] = 24'b000000000000100000100110 ; 
		block_ram[2087] = 24'b000001000000000010010000 ; 
		block_ram[2088] = 24'b000000000000100000101000 ; 
		block_ram[2089] = 24'b000000000000100000101001 ; 
		block_ram[2090] = 24'b000000000000100000101010 ; 
		block_ram[2091] = 24'b111000000000000000000000 ; 
		block_ram[2092] = 24'b000000000000100000101100 ; 
		block_ram[2093] = 24'b000000010000011000000000 ; 
		block_ram[2094] = 24'b000010000000000101000000 ; 
		block_ram[2095] = 24'b000000010000011000000010 ; 
		block_ram[2096] = 24'b000000000000100000110000 ; 
		block_ram[2097] = 24'b000000000000100000110001 ; 
		block_ram[2098] = 24'b000000000000100000110010 ; 
		block_ram[2099] = 24'b000001000000000010000100 ; 
		block_ram[2100] = 24'b000000000000100000110100 ; 
		block_ram[2101] = 24'b000001000000000010000010 ; 
		block_ram[2102] = 24'b000001000000000010000001 ; 
		block_ram[2103] = 24'b000001000000000010000000 ; 
		block_ram[2104] = 24'b000000000000100000111000 ; 
		block_ram[2105] = 24'b000110000100000000000000 ; 
		block_ram[2106] = 24'b000000000011001000000000 ; 
		block_ram[2107] = 24'b000000000011001000000001 ; 
		block_ram[2108] = 24'b010000101000000000000000 ; 
		block_ram[2109] = 24'b000000010000011000010000 ; 
		block_ram[2110] = 24'b000000000011001000000100 ; 
		block_ram[2111] = 24'b000001000000000010001000 ; 
		block_ram[2112] = 24'b000000000000100001000000 ; 
		block_ram[2113] = 24'b000000000000100001000001 ; 
		block_ram[2114] = 24'b000000000000100001000010 ; 
		block_ram[2115] = 24'b000000000000100001000011 ; 
		block_ram[2116] = 24'b000000000000100001000100 ; 
		block_ram[2117] = 24'b000000000000100001000101 ; 
		block_ram[2118] = 24'b000000000000100001000110 ; 
		block_ram[2119] = 24'b001000000001001000000000 ; 
		block_ram[2120] = 24'b000000000000100001001000 ; 
		block_ram[2121] = 24'b000000000000100001001001 ; 
		block_ram[2122] = 24'b000000000000100001001010 ; 
		block_ram[2123] = 24'b000000100000010000010000 ; 
		block_ram[2124] = 24'b000000000000100001001100 ; 
		block_ram[2125] = 24'b010001000100000000000000 ; 
		block_ram[2126] = 24'b000010000000000100100000 ; 
		block_ram[2127] = 24'b000000100000010000010100 ; 
		block_ram[2128] = 24'b000000000000100001010000 ; 
		block_ram[2129] = 24'b000000000000100001010001 ; 
		block_ram[2130] = 24'b000000000000100001010010 ; 
		block_ram[2131] = 24'b000000100000010000001000 ; 
		block_ram[2132] = 24'b000000000000100001010100 ; 
		block_ram[2133] = 24'b000010011000000000000000 ; 
		block_ram[2134] = 24'b110000000010000000000000 ; 
		block_ram[2135] = 24'b000000100000010000001100 ; 
		block_ram[2136] = 24'b000000000000100001011000 ; 
		block_ram[2137] = 24'b000000100000010000000010 ; 
		block_ram[2138] = 24'b000000100000010000000001 ; 
		block_ram[2139] = 24'b000000100000010000000000 ; 
		block_ram[2140] = 24'b000100000000001010000000 ; 
		block_ram[2141] = 24'b000000100000010000000110 ; 
		block_ram[2142] = 24'b000000100000010000000101 ; 
		block_ram[2143] = 24'b000000100000010000000100 ; 
		block_ram[2144] = 24'b000000000000100001100000 ; 
		block_ram[2145] = 24'b000000000000100001100001 ; 
		block_ram[2146] = 24'b000000000000100001100010 ; 
		block_ram[2147] = 24'b000000010110000000000000 ; 
		block_ram[2148] = 24'b000000000000100001100100 ; 
		block_ram[2149] = 24'b100100100000000000000000 ; 
		block_ram[2150] = 24'b000010000000000100001000 ; 
		block_ram[2151] = 24'b000000010110000000000100 ; 
		block_ram[2152] = 24'b000000000000100001101000 ; 
		block_ram[2153] = 24'b000000001001000010000000 ; 
		block_ram[2154] = 24'b000010000000000100000100 ; 
		block_ram[2155] = 24'b000000001001000010000010 ; 
		block_ram[2156] = 24'b000010000000000100000010 ; 
		block_ram[2157] = 24'b000000001001000010000100 ; 
		block_ram[2158] = 24'b000010000000000100000000 ; 
		block_ram[2159] = 24'b000010000000000100000001 ; 
		block_ram[2160] = 24'b000000000000100001110000 ; 
		block_ram[2161] = 24'b010000000000001100000000 ; 
		block_ram[2162] = 24'b001100001000000000000000 ; 
		block_ram[2163] = 24'b000000010110000000010000 ; 
		block_ram[2164] = 24'b000000000101010000000000 ; 
		block_ram[2165] = 24'b000000000101010000000001 ; 
		block_ram[2166] = 24'b000000000101010000000010 ; 
		block_ram[2167] = 24'b000001000000000011000000 ; 
		block_ram[2168] = 24'b100001010000000000000000 ; 
		block_ram[2169] = 24'b000000001001000010010000 ; 
		block_ram[2170] = 24'b000000000011001001000000 ; 
		block_ram[2171] = 24'b000000100000010000100000 ; 
		block_ram[2172] = 24'b000000000101010000001000 ; 
		block_ram[2173] = 24'b001000000010100000000000 ; 
		block_ram[2174] = 24'b000010000000000100010000 ; 
		block_ram[2175] = 24'b000000100000010000100100 ; 
		block_ram[2176] = 24'b000000000000100010000000 ; 
		block_ram[2177] = 24'b000000000000100010000001 ; 
		block_ram[2178] = 24'b000000000000100010000010 ; 
		block_ram[2179] = 24'b000000000000100010000011 ; 
		block_ram[2180] = 24'b000000000000100010000100 ; 
		block_ram[2181] = 24'b000000000000100010000101 ; 
		block_ram[2182] = 24'b000000000000100010000110 ; 
		block_ram[2183] = 24'b000001000000000000110000 ; 
		block_ram[2184] = 24'b000000000000100010001000 ; 
		block_ram[2185] = 24'b000000000000100010001001 ; 
		block_ram[2186] = 24'b000000000000100010001010 ; 
		block_ram[2187] = 24'b000000000100001100000000 ; 
		block_ram[2188] = 24'b000000000000100010001100 ; 
		block_ram[2189] = 24'b001010100000000000000000 ; 
		block_ram[2190] = 24'b010000000001010000000000 ; 
		block_ram[2191] = 24'b000000000100001100000100 ; 
		block_ram[2192] = 24'b000000000000100010010000 ; 
		block_ram[2193] = 24'b000000000000100010010001 ; 
		block_ram[2194] = 24'b000000000000100010010010 ; 
		block_ram[2195] = 24'b000001000000000000100100 ; 
		block_ram[2196] = 24'b000000000000100010010100 ; 
		block_ram[2197] = 24'b000001000000000000100010 ; 
		block_ram[2198] = 24'b000001000000000000100001 ; 
		block_ram[2199] = 24'b000001000000000000100000 ; 
		block_ram[2200] = 24'b000000000000100010011000 ; 
		block_ram[2201] = 24'b010000010010000000000000 ; 
		block_ram[2202] = 24'b100010001000000000000000 ; 
		block_ram[2203] = 24'b000000000100001100010000 ; 
		block_ram[2204] = 24'b000100000000001001000000 ; 
		block_ram[2205] = 24'b000000001100110000000000 ; 
		block_ram[2206] = 24'b000000100010100100000000 ; 
		block_ram[2207] = 24'b000001000000000000101000 ; 
		block_ram[2208] = 24'b000000000000100010100000 ; 
		block_ram[2209] = 24'b000000000000100010100001 ; 
		block_ram[2210] = 24'b000000000000100010100010 ; 
		block_ram[2211] = 24'b000001000000000000010100 ; 
		block_ram[2212] = 24'b000000000000100010100100 ; 
		block_ram[2213] = 24'b000001000000000000010010 ; 
		block_ram[2214] = 24'b000001000000000000010001 ; 
		block_ram[2215] = 24'b000001000000000000010000 ; 
		block_ram[2216] = 24'b000000000000100010101000 ; 
		block_ram[2217] = 24'b000000001001000001000000 ; 
		block_ram[2218] = 24'b000100110000000000000000 ; 
		block_ram[2219] = 24'b000000000100001100100000 ; 
		block_ram[2220] = 24'b100000000110000000000000 ; 
		block_ram[2221] = 24'b000000001001000001000100 ; 
		block_ram[2222] = 24'b000001000000000000011001 ; 
		block_ram[2223] = 24'b000001000000000000011000 ; 
		block_ram[2224] = 24'b000000000000100010110000 ; 
		block_ram[2225] = 24'b000001000000000000000110 ; 
		block_ram[2226] = 24'b000001000000000000000101 ; 
		block_ram[2227] = 24'b000001000000000000000100 ; 
		block_ram[2228] = 24'b000001000000000000000011 ; 
		block_ram[2229] = 24'b000001000000000000000010 ; 
		block_ram[2230] = 24'b000001000000000000000001 ; 
		block_ram[2231] = 24'b000001000000000000000000 ; 
		block_ram[2232] = 24'b001000000000010100000000 ; 
		block_ram[2233] = 24'b000000001001000001010000 ; 
		block_ram[2234] = 24'b000000000011001010000000 ; 
		block_ram[2235] = 24'b000001000000000000001100 ; 
		block_ram[2236] = 24'b000001000000000000001011 ; 
		block_ram[2237] = 24'b000001000000000000001010 ; 
		block_ram[2238] = 24'b000001000000000000001001 ; 
		block_ram[2239] = 24'b000001000000000000001000 ; 
		block_ram[2240] = 24'b000000000000100011000000 ; 
		block_ram[2241] = 24'b000000000000100011000001 ; 
		block_ram[2242] = 24'b000000000000100011000010 ; 
		block_ram[2243] = 24'b010110000000000000000000 ; 
		block_ram[2244] = 24'b000000000000100011000100 ; 
		block_ram[2245] = 24'b000000000010010100000000 ; 
		block_ram[2246] = 24'b000000101100000000000000 ; 
		block_ram[2247] = 24'b000000000010010100000010 ; 
		block_ram[2248] = 24'b000000000000100011001000 ; 
		block_ram[2249] = 24'b000000001001000000100000 ; 
		block_ram[2250] = 24'b001001000010000000000000 ; 
		block_ram[2251] = 24'b000000000100001101000000 ; 
		block_ram[2252] = 24'b000100000000001000010000 ; 
		block_ram[2253] = 24'b000000000010010100001000 ; 
		block_ram[2254] = 24'b000000101100000000001000 ; 
		block_ram[2255] = 24'b100000010000100000000000 ; 
		block_ram[2256] = 24'b000000000000100011010000 ; 
		block_ram[2257] = 24'b101000000100000000000000 ; 
		block_ram[2258] = 24'b000000010001000100000000 ; 
		block_ram[2259] = 24'b000000001010101000000000 ; 
		block_ram[2260] = 24'b000100000000001000001000 ; 
		block_ram[2261] = 24'b000000000010010100010000 ; 
		block_ram[2262] = 24'b000000010001000100000100 ; 
		block_ram[2263] = 24'b000001000000000001100000 ; 
		block_ram[2264] = 24'b000100000000001000000100 ; 
		block_ram[2265] = 24'b000000001001000000110000 ; 
		block_ram[2266] = 24'b000000010001000100001000 ; 
		block_ram[2267] = 24'b000000100000010010000000 ; 
		block_ram[2268] = 24'b000100000000001000000000 ; 
		block_ram[2269] = 24'b000100000000001000000001 ; 
		block_ram[2270] = 24'b000100000000001000000010 ; 
		block_ram[2271] = 24'b000000100000010010000100 ; 
		block_ram[2272] = 24'b000000000000100011100000 ; 
		block_ram[2273] = 24'b000000001001000000001000 ; 
		block_ram[2274] = 24'b100000000000011000000000 ; 
		block_ram[2275] = 24'b000000001001000000001010 ; 
		block_ram[2276] = 24'b011000010000000000000000 ; 
		block_ram[2277] = 24'b000000000010010100100000 ; 
		block_ram[2278] = 24'b000000101100000000100000 ; 
		block_ram[2279] = 24'b000001000000000001010000 ; 
		block_ram[2280] = 24'b000000001001000000000001 ; 
		block_ram[2281] = 24'b000000001001000000000000 ; 
		block_ram[2282] = 24'b000000001001000000000011 ; 
		block_ram[2283] = 24'b000000001001000000000010 ; 
		block_ram[2284] = 24'b000000001001000000000101 ; 
		block_ram[2285] = 24'b000000001001000000000100 ; 
		block_ram[2286] = 24'b000010000000000110000000 ; 
		block_ram[2287] = 24'b000000001001000000000110 ; 
		block_ram[2288] = 24'b000010100010000000000000 ; 
		block_ram[2289] = 24'b000000001001000000011000 ; 
		block_ram[2290] = 24'b000000010001000100100000 ; 
		block_ram[2291] = 24'b000001000000000001000100 ; 
		block_ram[2292] = 24'b000000000101010010000000 ; 
		block_ram[2293] = 24'b000001000000000001000010 ; 
		block_ram[2294] = 24'b000001000000000001000001 ; 
		block_ram[2295] = 24'b000001000000000001000000 ; 
		block_ram[2296] = 24'b000000001001000000010001 ; 
		block_ram[2297] = 24'b000000001001000000010000 ; 
		block_ram[2298] = 24'b010000000100100000000000 ; 
		block_ram[2299] = 24'b000000001001000000010010 ; 
		block_ram[2300] = 24'b000100000000001000100000 ; 
		block_ram[2301] = 24'b000000001001000000010100 ; 
		block_ram[2302] = 24'b000000011010010000000000 ; 
		block_ram[2303] = 24'b000001000000000001001000 ; 
		block_ram[2304] = 24'b000000000000100100000000 ; 
		block_ram[2305] = 24'b000000000000100100000001 ; 
		block_ram[2306] = 24'b000000000000100100000010 ; 
		block_ram[2307] = 24'b000000000000100100000011 ; 
		block_ram[2308] = 24'b000000000000100100000100 ; 
		block_ram[2309] = 24'b000000000000100100000101 ; 
		block_ram[2310] = 24'b000000000000100100000110 ; 
		block_ram[2311] = 24'b010000110000000000000000 ; 
		block_ram[2312] = 24'b000000000000100100001000 ; 
		block_ram[2313] = 24'b000000000000100100001001 ; 
		block_ram[2314] = 24'b000000000000100100001010 ; 
		block_ram[2315] = 24'b000000000100001010000000 ; 
		block_ram[2316] = 24'b000000000000100100001100 ; 
		block_ram[2317] = 24'b100000000001000000010000 ; 
		block_ram[2318] = 24'b000010000000000001100000 ; 
		block_ram[2319] = 24'b000000000100001010000100 ; 
		block_ram[2320] = 24'b000000000000100100010000 ; 
		block_ram[2321] = 24'b000000000000100100010001 ; 
		block_ram[2322] = 24'b000000000000100100010010 ; 
		block_ram[2323] = 24'b001010000010000000000000 ; 
		block_ram[2324] = 24'b000000000000100100010100 ; 
		block_ram[2325] = 24'b100000000001000000001000 ; 
		block_ram[2326] = 24'b000000001000011000000000 ; 
		block_ram[2327] = 24'b000000001000011000000001 ; 
		block_ram[2328] = 24'b000000000000100100011000 ; 
		block_ram[2329] = 24'b100000000001000000000100 ; 
		block_ram[2330] = 24'b010101000000000000000000 ; 
		block_ram[2331] = 24'b000000000100001010010000 ; 
		block_ram[2332] = 24'b100000000001000000000001 ; 
		block_ram[2333] = 24'b100000000001000000000000 ; 
		block_ram[2334] = 24'b000000001000011000001000 ; 
		block_ram[2335] = 24'b100000000001000000000010 ; 
		block_ram[2336] = 24'b000000000000100100100000 ; 
		block_ram[2337] = 24'b000000000000100100100001 ; 
		block_ram[2338] = 24'b000000000000100100100010 ; 
		block_ram[2339] = 24'b000100000001010000000000 ; 
		block_ram[2340] = 24'b000000000000100100100100 ; 
		block_ram[2341] = 24'b001000001100000000000000 ; 
		block_ram[2342] = 24'b000010000000000001001000 ; 
		block_ram[2343] = 24'b000001000000000110010000 ; 
		block_ram[2344] = 24'b000000000000100100101000 ; 
		block_ram[2345] = 24'b000001100010000000000000 ; 
		block_ram[2346] = 24'b000010000000000001000100 ; 
		block_ram[2347] = 24'b000000000100001010100000 ; 
		block_ram[2348] = 24'b000010000000000001000010 ; 
		block_ram[2349] = 24'b000000010000011100000000 ; 
		block_ram[2350] = 24'b000010000000000001000000 ; 
		block_ram[2351] = 24'b000010000000000001000001 ; 
		block_ram[2352] = 24'b000000000000100100110000 ; 
		block_ram[2353] = 24'b010000000000001001000000 ; 
		block_ram[2354] = 24'b100000100100000000000000 ; 
		block_ram[2355] = 24'b000000011000100000001000 ; 
		block_ram[2356] = 24'b000100010010000000000000 ; 
		block_ram[2357] = 24'b000001000000000110000010 ; 
		block_ram[2358] = 24'b000000001000011000100000 ; 
		block_ram[2359] = 24'b000001000000000110000000 ; 
		block_ram[2360] = 24'b001000000000010010000000 ; 
		block_ram[2361] = 24'b000000011000100000000010 ; 
		block_ram[2362] = 24'b000000000011001100000000 ; 
		block_ram[2363] = 24'b000000011000100000000000 ; 
		block_ram[2364] = 24'b000001000100101000000000 ; 
		block_ram[2365] = 24'b100000000001000000100000 ; 
		block_ram[2366] = 24'b000010000000000001010000 ; 
		block_ram[2367] = 24'b000000011000100000000100 ; 
		block_ram[2368] = 24'b000000000000100101000000 ; 
		block_ram[2369] = 24'b000000000000100101000001 ; 
		block_ram[2370] = 24'b000000000000100101000010 ; 
		block_ram[2371] = 24'b100001001000000000000000 ; 
		block_ram[2372] = 24'b000000000000100101000100 ; 
		block_ram[2373] = 24'b000000000010010010000000 ; 
		block_ram[2374] = 24'b000010000000000000101000 ; 
		block_ram[2375] = 24'b000000000010010010000010 ; 
		block_ram[2376] = 24'b000000000000100101001000 ; 
		block_ram[2377] = 24'b001100010000000000000000 ; 
		block_ram[2378] = 24'b000010000000000000100100 ; 
		block_ram[2379] = 24'b000000000100001011000000 ; 
		block_ram[2380] = 24'b000010000000000000100010 ; 
		block_ram[2381] = 24'b000000000010010010001000 ; 
		block_ram[2382] = 24'b000010000000000000100000 ; 
		block_ram[2383] = 24'b000010000000000000100001 ; 
		block_ram[2384] = 24'b000000000000100101010000 ; 
		block_ram[2385] = 24'b010000000000001000100000 ; 
		block_ram[2386] = 24'b000000010001000010000000 ; 
		block_ram[2387] = 24'b000000010001000010000001 ; 
		block_ram[2388] = 24'b001001100000000000000000 ; 
		block_ram[2389] = 24'b000000000010010010010000 ; 
		block_ram[2390] = 24'b000000001000011001000000 ; 
		block_ram[2391] = 24'b000100000100100000000000 ; 
		block_ram[2392] = 24'b000000001110000000000000 ; 
		block_ram[2393] = 24'b000000001110000000000001 ; 
		block_ram[2394] = 24'b000000001110000000000010 ; 
		block_ram[2395] = 24'b000000100000010100000000 ; 
		block_ram[2396] = 24'b000000001110000000000100 ; 
		block_ram[2397] = 24'b100000000001000001000000 ; 
		block_ram[2398] = 24'b000010000000000000110000 ; 
		block_ram[2399] = 24'b000000100000010100000100 ; 
		block_ram[2400] = 24'b000000000000100101100000 ; 
		block_ram[2401] = 24'b010000000000001000010000 ; 
		block_ram[2402] = 24'b000010000000000000001100 ; 
		block_ram[2403] = 24'b000000010110000100000000 ; 
		block_ram[2404] = 24'b000010000000000000001010 ; 
		block_ram[2405] = 24'b000000000010010010100000 ; 
		block_ram[2406] = 24'b000010000000000000001000 ; 
		block_ram[2407] = 24'b000010000000000000001001 ; 
		block_ram[2408] = 24'b000010000000000000000110 ; 
		block_ram[2409] = 24'b000000001001000110000000 ; 
		block_ram[2410] = 24'b000010000000000000000100 ; 
		block_ram[2411] = 24'b000010000000000000000101 ; 
		block_ram[2412] = 24'b000010000000000000000010 ; 
		block_ram[2413] = 24'b000010000000000000000011 ; 
		block_ram[2414] = 24'b000010000000000000000000 ; 
		block_ram[2415] = 24'b000010000000000000000001 ; 
		block_ram[2416] = 24'b010000000000001000000001 ; 
		block_ram[2417] = 24'b010000000000001000000000 ; 
		block_ram[2418] = 24'b000000010001000010100000 ; 
		block_ram[2419] = 24'b010000000000001000000010 ; 
		block_ram[2420] = 24'b000000000101010100000000 ; 
		block_ram[2421] = 24'b010000000000001000000100 ; 
		block_ram[2422] = 24'b000010000000000000011000 ; 
		block_ram[2423] = 24'b000000101011000000000000 ; 
		block_ram[2424] = 24'b000000001110000000100000 ; 
		block_ram[2425] = 24'b010000000000001000001000 ; 
		block_ram[2426] = 24'b000010000000000000010100 ; 
		block_ram[2427] = 24'b000000011000100001000000 ; 
		block_ram[2428] = 24'b000010000000000000010010 ; 
		block_ram[2429] = 24'b000000110100000010000000 ; 
		block_ram[2430] = 24'b000010000000000000010000 ; 
		block_ram[2431] = 24'b000010000000000000010001 ; 
		block_ram[2432] = 24'b000000000000100110000000 ; 
		block_ram[2433] = 24'b000000000000100110000001 ; 
		block_ram[2434] = 24'b000000000000100110000010 ; 
		block_ram[2435] = 24'b000000000100001000001000 ; 
		block_ram[2436] = 24'b000000000000100110000100 ; 
		block_ram[2437] = 24'b000000000010010001000000 ; 
		block_ram[2438] = 24'b101100000000000000000000 ; 
		block_ram[2439] = 24'b000000000010010001000010 ; 
		block_ram[2440] = 24'b000000000000100110001000 ; 
		block_ram[2441] = 24'b000000000100001000000010 ; 
		block_ram[2442] = 24'b000000000100001000000001 ; 
		block_ram[2443] = 24'b000000000100001000000000 ; 
		block_ram[2444] = 24'b000001011000000000000000 ; 
		block_ram[2445] = 24'b000000000010010001001000 ; 
		block_ram[2446] = 24'b000000000100001000000101 ; 
		block_ram[2447] = 24'b000000000100001000000100 ; 
		block_ram[2448] = 24'b000000000000100110010000 ; 
		block_ram[2449] = 24'b000100101000000000000000 ; 
		block_ram[2450] = 24'b000000010001000001000000 ; 
		block_ram[2451] = 24'b000000000100001000011000 ; 
		block_ram[2452] = 24'b010010000100000000000000 ; 
		block_ram[2453] = 24'b000000000010010001010000 ; 
		block_ram[2454] = 24'b000000001000011010000000 ; 
		block_ram[2455] = 24'b000001000000000100100000 ; 
		block_ram[2456] = 24'b001000000000010000100000 ; 
		block_ram[2457] = 24'b000000000100001000010010 ; 
		block_ram[2458] = 24'b000000000100001000010001 ; 
		block_ram[2459] = 24'b000000000100001000010000 ; 
		block_ram[2460] = 24'b000000100010100000000010 ; 
		block_ram[2461] = 24'b100000000001000010000000 ; 
		block_ram[2462] = 24'b000000100010100000000000 ; 
		block_ram[2463] = 24'b000000000100001000010100 ; 
		block_ram[2464] = 24'b000000000000100110100000 ; 
		block_ram[2465] = 24'b100010010000000000000000 ; 
		block_ram[2466] = 24'b010000001010000000000000 ; 
		block_ram[2467] = 24'b000000000100001000101000 ; 
		block_ram[2468] = 24'b000000100001001000000000 ; 
		block_ram[2469] = 24'b000000000010010001100000 ; 
		block_ram[2470] = 24'b000000010100110000000000 ; 
		block_ram[2471] = 24'b000001000000000100010000 ; 
		block_ram[2472] = 24'b001000000000010000010000 ; 
		block_ram[2473] = 24'b000000000100001000100010 ; 
		block_ram[2474] = 24'b000000000100001000100001 ; 
		block_ram[2475] = 24'b000000000100001000100000 ; 
		block_ram[2476] = 24'b000000100001001000001000 ; 
		block_ram[2477] = 24'b010100000000100000000000 ; 
		block_ram[2478] = 24'b000010000000000011000000 ; 
		block_ram[2479] = 24'b000000000100001000100100 ; 
		block_ram[2480] = 24'b001000000000010000001000 ; 
		block_ram[2481] = 24'b000000000111100000000000 ; 
		block_ram[2482] = 24'b000000010001000001100000 ; 
		block_ram[2483] = 24'b000001000000000100000100 ; 
		block_ram[2484] = 24'b000000100001001000010000 ; 
		block_ram[2485] = 24'b000001000000000100000010 ; 
		block_ram[2486] = 24'b000001000000000100000001 ; 
		block_ram[2487] = 24'b000001000000000100000000 ; 
		block_ram[2488] = 24'b001000000000010000000000 ; 
		block_ram[2489] = 24'b001000000000010000000001 ; 
		block_ram[2490] = 24'b001000000000010000000010 ; 
		block_ram[2491] = 24'b000000000100001000110000 ; 
		block_ram[2492] = 24'b001000000000010000000100 ; 
		block_ram[2493] = 24'b000000110100000001000000 ; 
		block_ram[2494] = 24'b000000100010100000100000 ; 
		block_ram[2495] = 24'b000001000000000100001000 ; 
		block_ram[2496] = 24'b000000000000100111000000 ; 
		block_ram[2497] = 24'b000000000010010000000100 ; 
		block_ram[2498] = 24'b000000010001000000010000 ; 
		block_ram[2499] = 24'b000000000010010000000110 ; 
		block_ram[2500] = 24'b000000000010010000000001 ; 
		block_ram[2501] = 24'b000000000010010000000000 ; 
		block_ram[2502] = 24'b000000000010010000000011 ; 
		block_ram[2503] = 24'b000000000010010000000010 ; 
		block_ram[2504] = 24'b110000100000000000000000 ; 
		block_ram[2505] = 24'b000000000010010000001100 ; 
		block_ram[2506] = 24'b000000000100001001000001 ; 
		block_ram[2507] = 24'b000000000100001001000000 ; 
		block_ram[2508] = 24'b000000000010010000001001 ; 
		block_ram[2509] = 24'b000000000010010000001000 ; 
		block_ram[2510] = 24'b000010000000000010100000 ; 
		block_ram[2511] = 24'b000000000010010000001010 ; 
		block_ram[2512] = 24'b000000010001000000000010 ; 
		block_ram[2513] = 24'b000000000010010000010100 ; 
		block_ram[2514] = 24'b000000010001000000000000 ; 
		block_ram[2515] = 24'b000000010001000000000001 ; 
		block_ram[2516] = 24'b000000000010010000010001 ; 
		block_ram[2517] = 24'b000000000010010000010000 ; 
		block_ram[2518] = 24'b000000010001000000000100 ; 
		block_ram[2519] = 24'b000000000010010000010010 ; 
		block_ram[2520] = 24'b000000001110000010000000 ; 
		block_ram[2521] = 24'b000011000000100000000000 ; 
		block_ram[2522] = 24'b000000010001000000001000 ; 
		block_ram[2523] = 24'b000000000100001001010000 ; 
		block_ram[2524] = 24'b000100000000001100000000 ; 
		block_ram[2525] = 24'b000000000010010000011000 ; 
		block_ram[2526] = 24'b000000010001000000001100 ; 
		block_ram[2527] = 24'b011000001000000000000000 ; 
		block_ram[2528] = 24'b000101000100000000000000 ; 
		block_ram[2529] = 24'b000000000010010000100100 ; 
		block_ram[2530] = 24'b000000010001000000110000 ; 
		block_ram[2531] = 24'b001000100000100000000000 ; 
		block_ram[2532] = 24'b000000000010010000100001 ; 
		block_ram[2533] = 24'b000000000010010000100000 ; 
		block_ram[2534] = 24'b000010000000000010001000 ; 
		block_ram[2535] = 24'b000000000010010000100010 ; 
		block_ram[2536] = 24'b000000001001000100000001 ; 
		block_ram[2537] = 24'b000000001001000100000000 ; 
		block_ram[2538] = 24'b000010000000000010000100 ; 
		block_ram[2539] = 24'b000000000100001001100000 ; 
		block_ram[2540] = 24'b000010000000000010000010 ; 
		block_ram[2541] = 24'b000000000010010000101000 ; 
		block_ram[2542] = 24'b000010000000000010000000 ; 
		block_ram[2543] = 24'b000010000000000010000001 ; 
		block_ram[2544] = 24'b000000010001000000100010 ; 
		block_ram[2545] = 24'b010000000000001010000000 ; 
		block_ram[2546] = 24'b000000010001000000100000 ; 
		block_ram[2547] = 24'b000000010001000000100001 ; 
		block_ram[2548] = 24'b100000001000100000000000 ; 
		block_ram[2549] = 24'b000000000010010000110000 ; 
		block_ram[2550] = 24'b000000010001000000100100 ; 
		block_ram[2551] = 24'b000001000000000101000000 ; 
		block_ram[2552] = 24'b001000000000010001000000 ; 
		block_ram[2553] = 24'b000000001001000100010000 ; 
		block_ram[2554] = 24'b000000010001000000101000 ; 
		block_ram[2555] = 24'b100100000010000000000000 ; 
		block_ram[2556] = 24'b000000110100000000000001 ; 
		block_ram[2557] = 24'b000000110100000000000000 ; 
		block_ram[2558] = 24'b000010000000000010010000 ; 
		block_ram[2559] = 24'b000000000001111000000000 ; 
		block_ram[2560] = 24'b000000000000101000000000 ; 
		block_ram[2561] = 24'b000000000000101000000001 ; 
		block_ram[2562] = 24'b000000000000101000000010 ; 
		block_ram[2563] = 24'b000000000000101000000011 ; 
		block_ram[2564] = 24'b000000000000101000000100 ; 
		block_ram[2565] = 24'b000000000000101000000101 ; 
		block_ram[2566] = 24'b000000000000101000000110 ; 
		block_ram[2567] = 24'b001000000001000001000000 ; 
		block_ram[2568] = 24'b000000000000101000001000 ; 
		block_ram[2569] = 24'b000000000000101000001001 ; 
		block_ram[2570] = 24'b000000000000101000001010 ; 
		block_ram[2571] = 24'b000000000100000110000000 ; 
		block_ram[2572] = 24'b000000000000101000001100 ; 
		block_ram[2573] = 24'b000000010000010000100000 ; 
		block_ram[2574] = 24'b100001100000000000000000 ; 
		block_ram[2575] = 24'b000000000100000110000100 ; 
		block_ram[2576] = 24'b000000000000101000010000 ; 
		block_ram[2577] = 24'b000000000000101000010001 ; 
		block_ram[2578] = 24'b000000000000101000010010 ; 
		block_ram[2579] = 24'b100100010000000000000000 ; 
		block_ram[2580] = 24'b000000000000101000010100 ; 
		block_ram[2581] = 24'b000000100110000000000000 ; 
		block_ram[2582] = 24'b000000001000010100000000 ; 
		block_ram[2583] = 24'b000000001000010100000001 ; 
		block_ram[2584] = 24'b000000000000101000011000 ; 
		block_ram[2585] = 24'b001001001000000000000000 ; 
		block_ram[2586] = 24'b000000000011000000100000 ; 
		block_ram[2587] = 24'b000000000011000000100001 ; 
		block_ram[2588] = 24'b000100000000000011000000 ; 
		block_ram[2589] = 24'b000000010000010000110000 ; 
		block_ram[2590] = 24'b000000000011000000100100 ; 
		block_ram[2591] = 24'b010010000000100000000000 ; 
		block_ram[2592] = 24'b000000000000101000100000 ; 
		block_ram[2593] = 24'b000000000000101000100001 ; 
		block_ram[2594] = 24'b000000000000101000100010 ; 
		block_ram[2595] = 24'b000010101000000000000000 ; 
		block_ram[2596] = 24'b000000000000101000100100 ; 
		block_ram[2597] = 24'b000000010000010000001000 ; 
		block_ram[2598] = 24'b010100000100000000000000 ; 
		block_ram[2599] = 24'b000000010000010000001010 ; 
		block_ram[2600] = 24'b000000000000101000101000 ; 
		block_ram[2601] = 24'b000000010000010000000100 ; 
		block_ram[2602] = 24'b000000000011000000010000 ; 
		block_ram[2603] = 24'b000000000011000000010001 ; 
		block_ram[2604] = 24'b000000010000010000000001 ; 
		block_ram[2605] = 24'b000000010000010000000000 ; 
		block_ram[2606] = 24'b000000000011000000010100 ; 
		block_ram[2607] = 24'b000000010000010000000010 ; 
		block_ram[2608] = 24'b000000000000101000110000 ; 
		block_ram[2609] = 24'b010000000000000101000000 ; 
		block_ram[2610] = 24'b000000000011000000001000 ; 
		block_ram[2611] = 24'b000000000011000000001001 ; 
		block_ram[2612] = 24'b101010000000000000000000 ; 
		block_ram[2613] = 24'b000000010000010000011000 ; 
		block_ram[2614] = 24'b000000000011000000001100 ; 
		block_ram[2615] = 24'b000001000000001010000000 ; 
		block_ram[2616] = 24'b000000000011000000000010 ; 
		block_ram[2617] = 24'b000000000011000000000011 ; 
		block_ram[2618] = 24'b000000000011000000000000 ; 
		block_ram[2619] = 24'b000000000011000000000001 ; 
		block_ram[2620] = 24'b000000000011000000000110 ; 
		block_ram[2621] = 24'b000000010000010000010000 ; 
		block_ram[2622] = 24'b000000000011000000000100 ; 
		block_ram[2623] = 24'b000000000011000000000101 ; 
		block_ram[2624] = 24'b000000000000101001000000 ; 
		block_ram[2625] = 24'b000000000000101001000001 ; 
		block_ram[2626] = 24'b000000000000101001000010 ; 
		block_ram[2627] = 24'b001000000001000000000100 ; 
		block_ram[2628] = 24'b000000000000101001000100 ; 
		block_ram[2629] = 24'b001000000001000000000010 ; 
		block_ram[2630] = 24'b001000000001000000000001 ; 
		block_ram[2631] = 24'b001000000001000000000000 ; 
		block_ram[2632] = 24'b000000000000101001001000 ; 
		block_ram[2633] = 24'b100010000010000000000000 ; 
		block_ram[2634] = 24'b010000011000000000000000 ; 
		block_ram[2635] = 24'b000000000100000111000000 ; 
		block_ram[2636] = 24'b000100000000000010010000 ; 
		block_ram[2637] = 24'b000000010000010001100000 ; 
		block_ram[2638] = 24'b000000000110110000000000 ; 
		block_ram[2639] = 24'b001000000001000000001000 ; 
		block_ram[2640] = 24'b000000000000101001010000 ; 
		block_ram[2641] = 24'b010000000000000100100000 ; 
		block_ram[2642] = 24'b000011000100000000000000 ; 
		block_ram[2643] = 24'b000000001010100010000000 ; 
		block_ram[2644] = 24'b000100000000000010001000 ; 
		block_ram[2645] = 24'b000000100110000001000000 ; 
		block_ram[2646] = 24'b000000001000010101000000 ; 
		block_ram[2647] = 24'b001000000001000000010000 ; 
		block_ram[2648] = 24'b000100000000000010000100 ; 
		block_ram[2649] = 24'b000000010101100000000000 ; 
		block_ram[2650] = 24'b000000000011000001100000 ; 
		block_ram[2651] = 24'b000000100000011000000000 ; 
		block_ram[2652] = 24'b000100000000000010000000 ; 
		block_ram[2653] = 24'b000100000000000010000001 ; 
		block_ram[2654] = 24'b000100000000000010000010 ; 
		block_ram[2655] = 24'b000000100000011000000100 ; 
		block_ram[2656] = 24'b000000000000101001100000 ; 
		block_ram[2657] = 24'b010000000000000100010000 ; 
		block_ram[2658] = 24'b100000000000010010000000 ; 
		block_ram[2659] = 24'b000000010110001000000000 ; 
		block_ram[2660] = 24'b000001001010000000000000 ; 
		block_ram[2661] = 24'b000000010000010001001000 ; 
		block_ram[2662] = 24'b000000110000100000010000 ; 
		block_ram[2663] = 24'b001000000001000000100000 ; 
		block_ram[2664] = 24'b001000100100000000000000 ; 
		block_ram[2665] = 24'b000000001001001010000000 ; 
		block_ram[2666] = 24'b000000000011000001010000 ; 
		block_ram[2667] = 24'b000101000000100000000000 ; 
		block_ram[2668] = 24'b000000010000010001000001 ; 
		block_ram[2669] = 24'b000000010000010001000000 ; 
		block_ram[2670] = 24'b000010000000001100000000 ; 
		block_ram[2671] = 24'b000000010000010001000010 ; 
		block_ram[2672] = 24'b010000000000000100000001 ; 
		block_ram[2673] = 24'b010000000000000100000000 ; 
		block_ram[2674] = 24'b000000000011000001001000 ; 
		block_ram[2675] = 24'b010000000000000100000010 ; 
		block_ram[2676] = 24'b000000000101011000000000 ; 
		block_ram[2677] = 24'b010000000000000100000100 ; 
		block_ram[2678] = 24'b000000110000100000000000 ; 
		block_ram[2679] = 24'b000000110000100000000001 ; 
		block_ram[2680] = 24'b000000000011000001000010 ; 
		block_ram[2681] = 24'b010000000000000100001000 ; 
		block_ram[2682] = 24'b000000000011000001000000 ; 
		block_ram[2683] = 24'b000000000011000001000001 ; 
		block_ram[2684] = 24'b000100000000000010100000 ; 
		block_ram[2685] = 24'b000000010000010001010000 ; 
		block_ram[2686] = 24'b000000000011000001000100 ; 
		block_ram[2687] = 24'b100000001100000000000000 ; 
		block_ram[2688] = 24'b000000000000101010000000 ; 
		block_ram[2689] = 24'b000000000000101010000001 ; 
		block_ram[2690] = 24'b000000000000101010000010 ; 
		block_ram[2691] = 24'b000000000100000100001000 ; 
		block_ram[2692] = 24'b000000000000101010000100 ; 
		block_ram[2693] = 24'b110000001000000000000000 ; 
		block_ram[2694] = 24'b000010010010000000000000 ; 
		block_ram[2695] = 24'b000000000100000100001100 ; 
		block_ram[2696] = 24'b000000000000101010001000 ; 
		block_ram[2697] = 24'b000000000100000100000010 ; 
		block_ram[2698] = 24'b000000000100000100000001 ; 
		block_ram[2699] = 24'b000000000100000100000000 ; 
		block_ram[2700] = 24'b000100000000000001010000 ; 
		block_ram[2701] = 24'b000000000100000100000110 ; 
		block_ram[2702] = 24'b000000000100000100000101 ; 
		block_ram[2703] = 24'b000000000100000100000100 ; 
		block_ram[2704] = 24'b000000000000101010010000 ; 
		block_ram[2705] = 24'b000010000001010000000000 ; 
		block_ram[2706] = 24'b011000100000000000000000 ; 
		block_ram[2707] = 24'b000000000100000100011000 ; 
		block_ram[2708] = 24'b000100000000000001001000 ; 
		block_ram[2709] = 24'b000000100110000010000000 ; 
		block_ram[2710] = 24'b000000001000010110000000 ; 
		block_ram[2711] = 24'b000001000000001000100000 ; 
		block_ram[2712] = 24'b000100000000000001000100 ; 
		block_ram[2713] = 24'b000000000100000100010010 ; 
		block_ram[2714] = 24'b000000000011000010100000 ; 
		block_ram[2715] = 24'b000000000100000100010000 ; 
		block_ram[2716] = 24'b000100000000000001000000 ; 
		block_ram[2717] = 24'b000100000000000001000001 ; 
		block_ram[2718] = 24'b000100000000000001000010 ; 
		block_ram[2719] = 24'b000000000100000100010100 ; 
		block_ram[2720] = 24'b000000000000101010100000 ; 
		block_ram[2721] = 24'b001100000010000000000000 ; 
		block_ram[2722] = 24'b100000000000010001000000 ; 
		block_ram[2723] = 24'b000000000100000100101000 ; 
		block_ram[2724] = 24'b000000100001000100000000 ; 
		block_ram[2725] = 24'b000000010000010010001000 ; 
		block_ram[2726] = 24'b000000100001000100000010 ; 
		block_ram[2727] = 24'b000001000000001000010000 ; 
		block_ram[2728] = 24'b010011000000000000000000 ; 
		block_ram[2729] = 24'b000000000100000100100010 ; 
		block_ram[2730] = 24'b000000000011000010010000 ; 
		block_ram[2731] = 24'b000000000100000100100000 ; 
		block_ram[2732] = 24'b000000010000010010000001 ; 
		block_ram[2733] = 24'b000000010000010010000000 ; 
		block_ram[2734] = 24'b001000001000100000000000 ; 
		block_ram[2735] = 24'b000000000100000100100100 ; 
		block_ram[2736] = 24'b000000011100000000000000 ; 
		block_ram[2737] = 24'b000000011100000000000001 ; 
		block_ram[2738] = 24'b000000000011000010001000 ; 
		block_ram[2739] = 24'b000001000000001000000100 ; 
		block_ram[2740] = 24'b000000011100000000000100 ; 
		block_ram[2741] = 24'b000001000000001000000010 ; 
		block_ram[2742] = 24'b000001000000001000000001 ; 
		block_ram[2743] = 24'b000001000000001000000000 ; 
		block_ram[2744] = 24'b000000000011000010000010 ; 
		block_ram[2745] = 24'b100000100000100000000000 ; 
		block_ram[2746] = 24'b000000000011000010000000 ; 
		block_ram[2747] = 24'b000000000011000010000001 ; 
		block_ram[2748] = 24'b000100000000000001100000 ; 
		block_ram[2749] = 24'b000000010000010010010000 ; 
		block_ram[2750] = 24'b000000000011000010000100 ; 
		block_ram[2751] = 24'b000001000000001000001000 ; 
		block_ram[2752] = 24'b000000000000101011000000 ; 
		block_ram[2753] = 24'b000001110000000000000000 ; 
		block_ram[2754] = 24'b100000000000010000100000 ; 
		block_ram[2755] = 24'b000000000100000101001000 ; 
		block_ram[2756] = 24'b000100000000000000011000 ; 
		block_ram[2757] = 24'b000000000010011100000000 ; 
		block_ram[2758] = 24'b000000101100001000000000 ; 
		block_ram[2759] = 24'b001000000001000010000000 ; 
		block_ram[2760] = 24'b000100000000000000010100 ; 
		block_ram[2761] = 24'b000000000100000101000010 ; 
		block_ram[2762] = 24'b000000000100000101000001 ; 
		block_ram[2763] = 24'b000000000100000101000000 ; 
		block_ram[2764] = 24'b000100000000000000010000 ; 
		block_ram[2765] = 24'b000100000000000000010001 ; 
		block_ram[2766] = 24'b000100000000000000010010 ; 
		block_ram[2767] = 24'b000000000100000101000100 ; 
		block_ram[2768] = 24'b000100000000000000001100 ; 
		block_ram[2769] = 24'b000000001010100000000010 ; 
		block_ram[2770] = 24'b000000001010100000000001 ; 
		block_ram[2771] = 24'b000000001010100000000000 ; 
		block_ram[2772] = 24'b000100000000000000001000 ; 
		block_ram[2773] = 24'b000100000000000000001001 ; 
		block_ram[2774] = 24'b000100000000000000001010 ; 
		block_ram[2775] = 24'b000000001010100000000100 ; 
		block_ram[2776] = 24'b000100000000000000000100 ; 
		block_ram[2777] = 24'b000100000000000000000101 ; 
		block_ram[2778] = 24'b000100000000000000000110 ; 
		block_ram[2779] = 24'b000000000100000101010000 ; 
		block_ram[2780] = 24'b000100000000000000000000 ; 
		block_ram[2781] = 24'b000100000000000000000001 ; 
		block_ram[2782] = 24'b000100000000000000000010 ; 
		block_ram[2783] = 24'b000100000000000000000011 ; 
		block_ram[2784] = 24'b100000000000010000000010 ; 
		block_ram[2785] = 24'b000000001001001000001000 ; 
		block_ram[2786] = 24'b100000000000010000000000 ; 
		block_ram[2787] = 24'b100000000000010000000001 ; 
		block_ram[2788] = 24'b000000100001000101000000 ; 
		block_ram[2789] = 24'b000010000100100000000000 ; 
		block_ram[2790] = 24'b100000000000010000000100 ; 
		block_ram[2791] = 24'b000001000000001001010000 ; 
		block_ram[2792] = 24'b000000001001001000000001 ; 
		block_ram[2793] = 24'b000000001001001000000000 ; 
		block_ram[2794] = 24'b100000000000010000001000 ; 
		block_ram[2795] = 24'b000000000100000101100000 ; 
		block_ram[2796] = 24'b000100000000000000110000 ; 
		block_ram[2797] = 24'b000000001001001000000100 ; 
		block_ram[2798] = 24'b000001010101000000000000 ; 
		block_ram[2799] = 24'b010000100010000000000000 ; 
		block_ram[2800] = 24'b000000011100000001000000 ; 
		block_ram[2801] = 24'b010000000000000110000000 ; 
		block_ram[2802] = 24'b100000000000010000010000 ; 
		block_ram[2803] = 24'b000000001010100000100000 ; 
		block_ram[2804] = 24'b000100000000000000101000 ; 
		block_ram[2805] = 24'b000001000000001001000010 ; 
		block_ram[2806] = 24'b000000110000100010000000 ; 
		block_ram[2807] = 24'b000001000000001001000000 ; 
		block_ram[2808] = 24'b000100000000000000100100 ; 
		block_ram[2809] = 24'b000000001001001000010000 ; 
		block_ram[2810] = 24'b000000000011000011000000 ; 
		block_ram[2811] = 24'b001010010000000000000000 ; 
		block_ram[2812] = 24'b000100000000000000100000 ; 
		block_ram[2813] = 24'b000100000000000000100001 ; 
		block_ram[2814] = 24'b000100000000000000100010 ; 
		block_ram[2815] = 24'b000000000001110100000000 ; 
		block_ram[2816] = 24'b000000000000101100000000 ; 
		block_ram[2817] = 24'b000000000000101100000001 ; 
		block_ram[2818] = 24'b000000000000101100000010 ; 
		block_ram[2819] = 24'b000000000100000010001000 ; 
		block_ram[2820] = 24'b000000000000101100000100 ; 
		block_ram[2821] = 24'b000111000000000000000000 ; 
		block_ram[2822] = 24'b000000001000010000010000 ; 
		block_ram[2823] = 24'b000000000100000010001100 ; 
		block_ram[2824] = 24'b000000000000101100001000 ; 
		block_ram[2825] = 24'b000000000100000010000010 ; 
		block_ram[2826] = 24'b000000000100000010000001 ; 
		block_ram[2827] = 24'b000000000100000010000000 ; 
		block_ram[2828] = 24'b011000000010000000000000 ; 
		block_ram[2829] = 24'b000000000100000010000110 ; 
		block_ram[2830] = 24'b000000000100000010000101 ; 
		block_ram[2831] = 24'b000000000100000010000100 ; 
		block_ram[2832] = 24'b000000000000101100010000 ; 
		block_ram[2833] = 24'b010000000000000001100000 ; 
		block_ram[2834] = 24'b000000001000010000000100 ; 
		block_ram[2835] = 24'b000000000100000010011000 ; 
		block_ram[2836] = 24'b000000001000010000000010 ; 
		block_ram[2837] = 24'b000000001000010000000011 ; 
		block_ram[2838] = 24'b000000001000010000000000 ; 
		block_ram[2839] = 24'b000000001000010000000001 ; 
		block_ram[2840] = 24'b000010110000000000000000 ; 
		block_ram[2841] = 24'b000000000100000010010010 ; 
		block_ram[2842] = 24'b000000000011000100100000 ; 
		block_ram[2843] = 24'b000000000100000010010000 ; 
		block_ram[2844] = 24'b000000001000010000001010 ; 
		block_ram[2845] = 24'b100000000001001000000000 ; 
		block_ram[2846] = 24'b000000001000010000001000 ; 
		block_ram[2847] = 24'b000000000100000010010100 ; 
		block_ram[2848] = 24'b000000000000101100100000 ; 
		block_ram[2849] = 24'b010000000000000001010000 ; 
		block_ram[2850] = 24'b001001010000000000000000 ; 
		block_ram[2851] = 24'b000000000100000010101000 ; 
		block_ram[2852] = 24'b000000100001000010000000 ; 
		block_ram[2853] = 24'b000000010000010100001000 ; 
		block_ram[2854] = 24'b000000001000010000110000 ; 
		block_ram[2855] = 24'b100000000010100000000000 ; 
		block_ram[2856] = 24'b100100001000000000000000 ; 
		block_ram[2857] = 24'b000000000100000010100010 ; 
		block_ram[2858] = 24'b000000000011000100010000 ; 
		block_ram[2859] = 24'b000000000100000010100000 ; 
		block_ram[2860] = 24'b000000010000010100000001 ; 
		block_ram[2861] = 24'b000000010000010100000000 ; 
		block_ram[2862] = 24'b000010000000001001000000 ; 
		block_ram[2863] = 24'b000000000100000010100100 ; 
		block_ram[2864] = 24'b010000000000000001000001 ; 
		block_ram[2865] = 24'b010000000000000001000000 ; 
		block_ram[2866] = 24'b000000000011000100001000 ; 
		block_ram[2867] = 24'b010000000000000001000010 ; 
		block_ram[2868] = 24'b000000001000010000100010 ; 
		block_ram[2869] = 24'b010000000000000001000100 ; 
		block_ram[2870] = 24'b000000001000010000100000 ; 
		block_ram[2871] = 24'b000000001000010000100001 ; 
		block_ram[2872] = 24'b000000000011000100000010 ; 
		block_ram[2873] = 24'b010000000000000001001000 ; 
		block_ram[2874] = 24'b000000000011000100000000 ; 
		block_ram[2875] = 24'b000000000011000100000001 ; 
		block_ram[2876] = 24'b000001000100100000000000 ; 
		block_ram[2877] = 24'b000000010000010100010000 ; 
		block_ram[2878] = 24'b000000000011000100000100 ; 
		block_ram[2879] = 24'b001100100000000000000000 ; 
		block_ram[2880] = 24'b000000000000101101000000 ; 
		block_ram[2881] = 24'b010000000000000000110000 ; 
		block_ram[2882] = 24'b000100100010000000000000 ; 
		block_ram[2883] = 24'b000000000100000011001000 ; 
		block_ram[2884] = 24'b100000010100000000000000 ; 
		block_ram[2885] = 24'b000000000010011010000000 ; 
		block_ram[2886] = 24'b000000001000010001010000 ; 
		block_ram[2887] = 24'b001000000001000100000000 ; 
		block_ram[2888] = 24'b000001000001010000000000 ; 
		block_ram[2889] = 24'b000000000100000011000010 ; 
		block_ram[2890] = 24'b000000000100000011000001 ; 
		block_ram[2891] = 24'b000000000100000011000000 ; 
		block_ram[2892] = 24'b000000101000100000000001 ; 
		block_ram[2893] = 24'b000000101000100000000000 ; 
		block_ram[2894] = 24'b000010000000001000100000 ; 
		block_ram[2895] = 24'b000000000100000011000100 ; 
		block_ram[2896] = 24'b010000000000000000100001 ; 
		block_ram[2897] = 24'b010000000000000000100000 ; 
		block_ram[2898] = 24'b000000001000010001000100 ; 
		block_ram[2899] = 24'b010000000000000000100010 ; 
		block_ram[2900] = 24'b000000001000010001000010 ; 
		block_ram[2901] = 24'b010000000000000000100100 ; 
		block_ram[2902] = 24'b000000001000010001000000 ; 
		block_ram[2903] = 24'b000000001000010001000001 ; 
		block_ram[2904] = 24'b000000001110001000000000 ; 
		block_ram[2905] = 24'b010000000000000000101000 ; 
		block_ram[2906] = 24'b101000000000100000000000 ; 
		block_ram[2907] = 24'b000000000100000011010000 ; 
		block_ram[2908] = 24'b000100000000000110000000 ; 
		block_ram[2909] = 24'b000000101000100000010000 ; 
		block_ram[2910] = 24'b000000001000010001001000 ; 
		block_ram[2911] = 24'b000001010010000000000000 ; 
		block_ram[2912] = 24'b010000000000000000010001 ; 
		block_ram[2913] = 24'b010000000000000000010000 ; 
		block_ram[2914] = 24'b000000001101100000000000 ; 
		block_ram[2915] = 24'b010000000000000000010010 ; 
		block_ram[2916] = 24'b000000100001000011000000 ; 
		block_ram[2917] = 24'b010000000000000000010100 ; 
		block_ram[2918] = 24'b000010000000001000001000 ; 
		block_ram[2919] = 24'b000001100100010000000000 ; 
		block_ram[2920] = 24'b000000010010100010000000 ; 
		block_ram[2921] = 24'b010000000000000000011000 ; 
		block_ram[2922] = 24'b000010000000001000000100 ; 
		block_ram[2923] = 24'b000000000100000011100000 ; 
		block_ram[2924] = 24'b000010000000001000000010 ; 
		block_ram[2925] = 24'b000000010000010101000000 ; 
		block_ram[2926] = 24'b000010000000001000000000 ; 
		block_ram[2927] = 24'b000010000000001000000001 ; 
		block_ram[2928] = 24'b010000000000000000000001 ; 
		block_ram[2929] = 24'b010000000000000000000000 ; 
		block_ram[2930] = 24'b010000000000000000000011 ; 
		block_ram[2931] = 24'b010000000000000000000010 ; 
		block_ram[2932] = 24'b010000000000000000000101 ; 
		block_ram[2933] = 24'b010000000000000000000100 ; 
		block_ram[2934] = 24'b000000001000010001100000 ; 
		block_ram[2935] = 24'b010000000000000000000110 ; 
		block_ram[2936] = 24'b010000000000000000001001 ; 
		block_ram[2937] = 24'b010000000000000000001000 ; 
		block_ram[2938] = 24'b000000000011000101000000 ; 
		block_ram[2939] = 24'b010000000000000000001010 ; 
		block_ram[2940] = 24'b000001000100100001000000 ; 
		block_ram[2941] = 24'b010000000000000000001100 ; 
		block_ram[2942] = 24'b000010000000001000010000 ; 
		block_ram[2943] = 24'b000000000001110010000000 ; 
		block_ram[2944] = 24'b000000000000101110000000 ; 
		block_ram[2945] = 24'b000000000100000000001010 ; 
		block_ram[2946] = 24'b000000000100000000001001 ; 
		block_ram[2947] = 24'b000000000100000000001000 ; 
		block_ram[2948] = 24'b000000100001000000100000 ; 
		block_ram[2949] = 24'b000000000010011001000000 ; 
		block_ram[2950] = 24'b000000000100000000001101 ; 
		block_ram[2951] = 24'b000000000100000000001100 ; 
		block_ram[2952] = 24'b000000000100000000000011 ; 
		block_ram[2953] = 24'b000000000100000000000010 ; 
		block_ram[2954] = 24'b000000000100000000000001 ; 
		block_ram[2955] = 24'b000000000100000000000000 ; 
		block_ram[2956] = 24'b000000000100000000000111 ; 
		block_ram[2957] = 24'b000000000100000000000110 ; 
		block_ram[2958] = 24'b000000000100000000000101 ; 
		block_ram[2959] = 24'b000000000100000000000100 ; 
		block_ram[2960] = 24'b100001000010000000000000 ; 
		block_ram[2961] = 24'b000000000100000000011010 ; 
		block_ram[2962] = 24'b000000000100000000011001 ; 
		block_ram[2963] = 24'b000000000100000000011000 ; 
		block_ram[2964] = 24'b000000001000010010000010 ; 
		block_ram[2965] = 24'b001000010000100000000000 ; 
		block_ram[2966] = 24'b000000001000010010000000 ; 
		block_ram[2967] = 24'b000000000100000000011100 ; 
		block_ram[2968] = 24'b000000000100000000010011 ; 
		block_ram[2969] = 24'b000000000100000000010010 ; 
		block_ram[2970] = 24'b000000000100000000010001 ; 
		block_ram[2971] = 24'b000000000100000000010000 ; 
		block_ram[2972] = 24'b000100000000000101000000 ; 
		block_ram[2973] = 24'b000000000100000000010110 ; 
		block_ram[2974] = 24'b000000000100000000010101 ; 
		block_ram[2975] = 24'b000000000100000000010100 ; 
		block_ram[2976] = 24'b000000100001000000000100 ; 
		block_ram[2977] = 24'b000000000100000000101010 ; 
		block_ram[2978] = 24'b000000000100000000101001 ; 
		block_ram[2979] = 24'b000000000100000000101000 ; 
		block_ram[2980] = 24'b000000100001000000000000 ; 
		block_ram[2981] = 24'b000000100001000000000001 ; 
		block_ram[2982] = 24'b000000100001000000000010 ; 
		block_ram[2983] = 24'b000000000100000000101100 ; 
		block_ram[2984] = 24'b000000000100000000100011 ; 
		block_ram[2985] = 24'b000000000100000000100010 ; 
		block_ram[2986] = 24'b000000000100000000100001 ; 
		block_ram[2987] = 24'b000000000100000000100000 ; 
		block_ram[2988] = 24'b000000100001000000001000 ; 
		block_ram[2989] = 24'b000000000100000000100110 ; 
		block_ram[2990] = 24'b000000000100000000100101 ; 
		block_ram[2991] = 24'b000000000100000000100100 ; 
		block_ram[2992] = 24'b000000011100000100000000 ; 
		block_ram[2993] = 24'b010000000000000011000000 ; 
		block_ram[2994] = 24'b000110000000100000000000 ; 
		block_ram[2995] = 24'b000000000100000000111000 ; 
		block_ram[2996] = 24'b000000100001000000010000 ; 
		block_ram[2997] = 24'b000000100001000000010001 ; 
		block_ram[2998] = 24'b000000001000010010100000 ; 
		block_ram[2999] = 24'b000001000000001100000000 ; 
		block_ram[3000] = 24'b001000000000011000000000 ; 
		block_ram[3001] = 24'b000000000100000000110010 ; 
		block_ram[3002] = 24'b000000000011000110000000 ; 
		block_ram[3003] = 24'b000000000100000000110000 ; 
		block_ram[3004] = 24'b000000100001000000011000 ; 
		block_ram[3005] = 24'b000010001010000000000000 ; 
		block_ram[3006] = 24'b110000010000000000000000 ; 
		block_ram[3007] = 24'b000000000001110001000000 ; 
		block_ram[3008] = 24'b001010001000000000000000 ; 
		block_ram[3009] = 24'b000000000010011000000100 ; 
		block_ram[3010] = 24'b000000000100000001001001 ; 
		block_ram[3011] = 24'b000000000100000001001000 ; 
		block_ram[3012] = 24'b000000000010011000000001 ; 
		block_ram[3013] = 24'b000000000010011000000000 ; 
		block_ram[3014] = 24'b010001000000100000000000 ; 
		block_ram[3015] = 24'b000000000010011000000010 ; 
		block_ram[3016] = 24'b000000000100000001000011 ; 
		block_ram[3017] = 24'b000000000100000001000010 ; 
		block_ram[3018] = 24'b000000000100000001000001 ; 
		block_ram[3019] = 24'b000000000100000001000000 ; 
		block_ram[3020] = 24'b000100000000000100010000 ; 
		block_ram[3021] = 24'b000000000010011000001000 ; 
		block_ram[3022] = 24'b000000000100000001000101 ; 
		block_ram[3023] = 24'b000000000100000001000100 ; 
		block_ram[3024] = 24'b000000010001001000000010 ; 
		block_ram[3025] = 24'b010000000000000010100000 ; 
		block_ram[3026] = 24'b000000010001001000000000 ; 
		block_ram[3027] = 24'b000000000100000001011000 ; 
		block_ram[3028] = 24'b000100000000000100001000 ; 
		block_ram[3029] = 24'b000000000010011000010000 ; 
		block_ram[3030] = 24'b000000001000010011000000 ; 
		block_ram[3031] = 24'b100010100000000000000000 ; 
		block_ram[3032] = 24'b000100000000000100000100 ; 
		block_ram[3033] = 24'b000000000100000001010010 ; 
		block_ram[3034] = 24'b000000000100000001010001 ; 
		block_ram[3035] = 24'b000000000100000001010000 ; 
		block_ram[3036] = 24'b000100000000000100000000 ; 
		block_ram[3037] = 24'b000100000000000100000001 ; 
		block_ram[3038] = 24'b000100000000000100000010 ; 
		block_ram[3039] = 24'b000000000001110000100000 ; 
		block_ram[3040] = 24'b000000010010100000001000 ; 
		block_ram[3041] = 24'b010000000000000010010000 ; 
		block_ram[3042] = 24'b100000000000010100000000 ; 
		block_ram[3043] = 24'b000000000100000001101000 ; 
		block_ram[3044] = 24'b000000100001000001000000 ; 
		block_ram[3045] = 24'b000000000010011000100000 ; 
		block_ram[3046] = 24'b000000100001000001000010 ; 
		block_ram[3047] = 24'b000100011000000000000000 ; 
		block_ram[3048] = 24'b000000010010100000000000 ; 
		block_ram[3049] = 24'b000000000100000001100010 ; 
		block_ram[3050] = 24'b000000000100000001100001 ; 
		block_ram[3051] = 24'b000000000100000001100000 ; 
		block_ram[3052] = 24'b000000010010100000000100 ; 
		block_ram[3053] = 24'b101001000000000000000000 ; 
		block_ram[3054] = 24'b000010000000001010000000 ; 
		block_ram[3055] = 24'b000000000001110000010000 ; 
		block_ram[3056] = 24'b010000000000000010000001 ; 
		block_ram[3057] = 24'b010000000000000010000000 ; 
		block_ram[3058] = 24'b000000010001001000100000 ; 
		block_ram[3059] = 24'b010000000000000010000010 ; 
		block_ram[3060] = 24'b000000100001000001010000 ; 
		block_ram[3061] = 24'b010000000000000010000100 ; 
		block_ram[3062] = 24'b001000000110000000000000 ; 
		block_ram[3063] = 24'b000000000001110000001000 ; 
		block_ram[3064] = 24'b000000010010100000010000 ; 
		block_ram[3065] = 24'b010000000000000010001000 ; 
		block_ram[3066] = 24'b000001101000000000000000 ; 
		block_ram[3067] = 24'b000000000001110000000100 ; 
		block_ram[3068] = 24'b000100000000000100100000 ; 
		block_ram[3069] = 24'b000000000001110000000010 ; 
		block_ram[3070] = 24'b000000000001110000000001 ; 
		block_ram[3071] = 24'b000000000001110000000000 ; 
		block_ram[3072] = 24'b000000000000110000000000 ; 
		block_ram[3073] = 24'b000000000000110000000001 ; 
		block_ram[3074] = 24'b000000000000110000000010 ; 
		block_ram[3075] = 24'b000000000000110000000011 ; 
		block_ram[3076] = 24'b000000000000110000000100 ; 
		block_ram[3077] = 24'b000000000000110000000101 ; 
		block_ram[3078] = 24'b000000000000110000000110 ; 
		block_ram[3079] = 24'b100010000100000000000000 ; 
		block_ram[3080] = 24'b000000000000110000001000 ; 
		block_ram[3081] = 24'b000000000000110000001001 ; 
		block_ram[3082] = 24'b000000000000110000001010 ; 
		block_ram[3083] = 24'b000000100000000001010000 ; 
		block_ram[3084] = 24'b000000000000110000001100 ; 
		block_ram[3085] = 24'b000000010000001000100000 ; 
		block_ram[3086] = 24'b010000000001000010000000 ; 
		block_ram[3087] = 24'b000000010000001000100010 ; 
		block_ram[3088] = 24'b000000000000110000010000 ; 
		block_ram[3089] = 24'b000000000000110000010001 ; 
		block_ram[3090] = 24'b000000000000110000010010 ; 
		block_ram[3091] = 24'b000000100000000001001000 ; 
		block_ram[3092] = 24'b000000000000110000010100 ; 
		block_ram[3093] = 24'b011100000000000000000000 ; 
		block_ram[3094] = 24'b000000001000001100000000 ; 
		block_ram[3095] = 24'b000000001000001100000001 ; 
		block_ram[3096] = 24'b000000000000110000011000 ; 
		block_ram[3097] = 24'b000000100000000001000010 ; 
		block_ram[3098] = 24'b000000100000000001000001 ; 
		block_ram[3099] = 24'b000000100000000001000000 ; 
		block_ram[3100] = 24'b000011000010000000000000 ; 
		block_ram[3101] = 24'b000000001100100010000000 ; 
		block_ram[3102] = 24'b000000001000001100001000 ; 
		block_ram[3103] = 24'b000000100000000001000100 ; 
		block_ram[3104] = 24'b000000000000110000100000 ; 
		block_ram[3105] = 24'b000000000000110000100001 ; 
		block_ram[3106] = 24'b000000000000110000100010 ; 
		block_ram[3107] = 24'b000100000001000100000000 ; 
		block_ram[3108] = 24'b000000000000110000100100 ; 
		block_ram[3109] = 24'b000000010000001000001000 ; 
		block_ram[3110] = 24'b001000100010000000000000 ; 
		block_ram[3111] = 24'b000000010000001000001010 ; 
		block_ram[3112] = 24'b000000000000110000101000 ; 
		block_ram[3113] = 24'b000000010000001000000100 ; 
		block_ram[3114] = 24'b000001001100000000000000 ; 
		block_ram[3115] = 24'b000000010000001000000110 ; 
		block_ram[3116] = 24'b000000010000001000000001 ; 
		block_ram[3117] = 24'b000000010000001000000000 ; 
		block_ram[3118] = 24'b000000010000001000000011 ; 
		block_ram[3119] = 24'b000000010000001000000010 ; 
		block_ram[3120] = 24'b000000000000110000110000 ; 
		block_ram[3121] = 24'b100000001010000000000000 ; 
		block_ram[3122] = 24'b010010010000000000000000 ; 
		block_ram[3123] = 24'b000000100000000001101000 ; 
		block_ram[3124] = 24'b000000000101000001000000 ; 
		block_ram[3125] = 24'b000000000101000001000001 ; 
		block_ram[3126] = 24'b000000000101000001000010 ; 
		block_ram[3127] = 24'b000001000000010010000000 ; 
		block_ram[3128] = 24'b001000000000000110000000 ; 
		block_ram[3129] = 24'b000000010000001000010100 ; 
		block_ram[3130] = 24'b000000000011011000000000 ; 
		block_ram[3131] = 24'b000000100000000001100000 ; 
		block_ram[3132] = 24'b000000000101000001001000 ; 
		block_ram[3133] = 24'b000000010000001000010000 ; 
		block_ram[3134] = 24'b100100000000100000000000 ; 
		block_ram[3135] = 24'b000000010000001000010010 ; 
		block_ram[3136] = 24'b000000000000110001000000 ; 
		block_ram[3137] = 24'b000000000000110001000001 ; 
		block_ram[3138] = 24'b000000000000110001000010 ; 
		block_ram[3139] = 24'b000000100000000000011000 ; 
		block_ram[3140] = 24'b000000000000110001000100 ; 
		block_ram[3141] = 24'b000000000010000110000000 ; 
		block_ram[3142] = 24'b000101010000000000000000 ; 
		block_ram[3143] = 24'b000000000010000110000010 ; 
		block_ram[3144] = 24'b000000000000110001001000 ; 
		block_ram[3145] = 24'b000000100000000000010010 ; 
		block_ram[3146] = 24'b000000100000000000010001 ; 
		block_ram[3147] = 24'b000000100000000000010000 ; 
		block_ram[3148] = 24'b101000001000000000000000 ; 
		block_ram[3149] = 24'b000000000010000110001000 ; 
		block_ram[3150] = 24'b000000000110101000000000 ; 
		block_ram[3151] = 24'b000000100000000000010100 ; 
		block_ram[3152] = 24'b000000000000110001010000 ; 
		block_ram[3153] = 24'b000000100000000000001010 ; 
		block_ram[3154] = 24'b000000100000000000001001 ; 
		block_ram[3155] = 24'b000000100000000000001000 ; 
		block_ram[3156] = 24'b000000000101000000100000 ; 
		block_ram[3157] = 24'b000000000010000110010000 ; 
		block_ram[3158] = 24'b000000000101000000100010 ; 
		block_ram[3159] = 24'b000000100000000000001100 ; 
		block_ram[3160] = 24'b000000100000000000000011 ; 
		block_ram[3161] = 24'b000000100000000000000010 ; 
		block_ram[3162] = 24'b000000100000000000000001 ; 
		block_ram[3163] = 24'b000000100000000000000000 ; 
		block_ram[3164] = 24'b000000000101000000101000 ; 
		block_ram[3165] = 24'b000000100000000000000110 ; 
		block_ram[3166] = 24'b000000100000000000000101 ; 
		block_ram[3167] = 24'b000000100000000000000100 ; 
		block_ram[3168] = 24'b000000000000110001100000 ; 
		block_ram[3169] = 24'b001011000000000000000000 ; 
		block_ram[3170] = 24'b100000000000001010000000 ; 
		block_ram[3171] = 24'b000000010110010000000000 ; 
		block_ram[3172] = 24'b000000000101000000010000 ; 
		block_ram[3173] = 24'b000000000010000110100000 ; 
		block_ram[3174] = 24'b000000000101000000010010 ; 
		block_ram[3175] = 24'b010000001000100000000000 ; 
		block_ram[3176] = 24'b010100000010000000000000 ; 
		block_ram[3177] = 24'b000000001001010010000000 ; 
		block_ram[3178] = 24'b000000100000000000110001 ; 
		block_ram[3179] = 24'b000000100000000000110000 ; 
		block_ram[3180] = 24'b000000000101000000011000 ; 
		block_ram[3181] = 24'b000000010000001001000000 ; 
		block_ram[3182] = 24'b000010000000010100000000 ; 
		block_ram[3183] = 24'b000000010000001001000010 ; 
		block_ram[3184] = 24'b000000000101000000000100 ; 
		block_ram[3185] = 24'b000000000101000000000101 ; 
		block_ram[3186] = 24'b000000000101000000000110 ; 
		block_ram[3187] = 24'b000000100000000000101000 ; 
		block_ram[3188] = 24'b000000000101000000000000 ; 
		block_ram[3189] = 24'b000000000101000000000001 ; 
		block_ram[3190] = 24'b000000000101000000000010 ; 
		block_ram[3191] = 24'b000000000101000000000011 ; 
		block_ram[3192] = 24'b000000000101000000001100 ; 
		block_ram[3193] = 24'b000000100000000000100010 ; 
		block_ram[3194] = 24'b000000100000000000100001 ; 
		block_ram[3195] = 24'b000000100000000000100000 ; 
		block_ram[3196] = 24'b000000000101000000001000 ; 
		block_ram[3197] = 24'b000000000101000000001001 ; 
		block_ram[3198] = 24'b000000000101000000001010 ; 
		block_ram[3199] = 24'b000000100000000000100100 ; 
		block_ram[3200] = 24'b000000000000110010000000 ; 
		block_ram[3201] = 24'b000000000000110010000001 ; 
		block_ram[3202] = 24'b000000000000110010000010 ; 
		block_ram[3203] = 24'b001000011000000000000000 ; 
		block_ram[3204] = 24'b000000000000110010000100 ; 
		block_ram[3205] = 24'b000000000010000101000000 ; 
		block_ram[3206] = 24'b010000000001000000001000 ; 
		block_ram[3207] = 24'b000000000010000101000010 ; 
		block_ram[3208] = 24'b000000000000110010001000 ; 
		block_ram[3209] = 24'b100101000000000000000000 ; 
		block_ram[3210] = 24'b010000000001000000000100 ; 
		block_ram[3211] = 24'b000000000100011100000000 ; 
		block_ram[3212] = 24'b010000000001000000000010 ; 
		block_ram[3213] = 24'b000000000010000101001000 ; 
		block_ram[3214] = 24'b010000000001000000000000 ; 
		block_ram[3215] = 24'b010000000001000000000001 ; 
		block_ram[3216] = 24'b000000000000110010010000 ; 
		block_ram[3217] = 24'b000010000001001000000000 ; 
		block_ram[3218] = 24'b000100000110000000000000 ; 
		block_ram[3219] = 24'b000000100000000011001000 ; 
		block_ram[3220] = 24'b100000110000000000000000 ; 
		block_ram[3221] = 24'b000000000010000101010000 ; 
		block_ram[3222] = 24'b000000001000001110000000 ; 
		block_ram[3223] = 24'b000001000000010000100000 ; 
		block_ram[3224] = 24'b001000000000000100100000 ; 
		block_ram[3225] = 24'b000000001100100000000100 ; 
		block_ram[3226] = 24'b000000100000000011000001 ; 
		block_ram[3227] = 24'b000000100000000011000000 ; 
		block_ram[3228] = 24'b000000001100100000000001 ; 
		block_ram[3229] = 24'b000000001100100000000000 ; 
		block_ram[3230] = 24'b010000000001000000010000 ; 
		block_ram[3231] = 24'b000000001100100000000010 ; 
		block_ram[3232] = 24'b000000000000110010100000 ; 
		block_ram[3233] = 24'b010000100100000000000000 ; 
		block_ram[3234] = 24'b100000000000001001000000 ; 
		block_ram[3235] = 24'b000001000000010000010100 ; 
		block_ram[3236] = 24'b000110001000000000000000 ; 
		block_ram[3237] = 24'b000000000010000101100000 ; 
		block_ram[3238] = 24'b000000010100100100000000 ; 
		block_ram[3239] = 24'b000001000000010000010000 ; 
		block_ram[3240] = 24'b001000000000000100010000 ; 
		block_ram[3241] = 24'b000000001001010001000000 ; 
		block_ram[3242] = 24'b000001001100000010000000 ; 
		block_ram[3243] = 24'b000010000010100000000000 ; 
		block_ram[3244] = 24'b000000010000001010000001 ; 
		block_ram[3245] = 24'b000000010000001010000000 ; 
		block_ram[3246] = 24'b010000000001000000100000 ; 
		block_ram[3247] = 24'b000000010000001010000010 ; 
		block_ram[3248] = 24'b001000000000000100001000 ; 
		block_ram[3249] = 24'b000001000000010000000110 ; 
		block_ram[3250] = 24'b000000101001100000000000 ; 
		block_ram[3251] = 24'b000001000000010000000100 ; 
		block_ram[3252] = 24'b000000000101000011000000 ; 
		block_ram[3253] = 24'b000001000000010000000010 ; 
		block_ram[3254] = 24'b000001000000010000000001 ; 
		block_ram[3255] = 24'b000001000000010000000000 ; 
		block_ram[3256] = 24'b001000000000000100000000 ; 
		block_ram[3257] = 24'b001000000000000100000001 ; 
		block_ram[3258] = 24'b001000000000000100000010 ; 
		block_ram[3259] = 24'b000000100000000011100000 ; 
		block_ram[3260] = 24'b001000000000000100000100 ; 
		block_ram[3261] = 24'b000000001100100000100000 ; 
		block_ram[3262] = 24'b000000011010000001000000 ; 
		block_ram[3263] = 24'b000001000000010000001000 ; 
		block_ram[3264] = 24'b000000000000110011000000 ; 
		block_ram[3265] = 24'b000000000010000100000100 ; 
		block_ram[3266] = 24'b100000000000001000100000 ; 
		block_ram[3267] = 24'b000000000010000100000110 ; 
		block_ram[3268] = 24'b000000000010000100000001 ; 
		block_ram[3269] = 24'b000000000010000100000000 ; 
		block_ram[3270] = 24'b000000000010000100000011 ; 
		block_ram[3271] = 24'b000000000010000100000010 ; 
		block_ram[3272] = 24'b000010010100000000000000 ; 
		block_ram[3273] = 24'b000000000010000100001100 ; 
		block_ram[3274] = 24'b000000100000000010010001 ; 
		block_ram[3275] = 24'b000000100000000010010000 ; 
		block_ram[3276] = 24'b000000000010000100001001 ; 
		block_ram[3277] = 24'b000000000010000100001000 ; 
		block_ram[3278] = 24'b010000000001000001000000 ; 
		block_ram[3279] = 24'b000000000010000100001010 ; 
		block_ram[3280] = 24'b010001001000000000000000 ; 
		block_ram[3281] = 24'b000000000010000100010100 ; 
		block_ram[3282] = 24'b000000010001010100000000 ; 
		block_ram[3283] = 24'b000000100000000010001000 ; 
		block_ram[3284] = 24'b000000000010000100010001 ; 
		block_ram[3285] = 24'b000000000010000100010000 ; 
		block_ram[3286] = 24'b001010000000100000000000 ; 
		block_ram[3287] = 24'b000000000010000100010010 ; 
		block_ram[3288] = 24'b000000100000000010000011 ; 
		block_ram[3289] = 24'b000000100000000010000010 ; 
		block_ram[3290] = 24'b000000100000000010000001 ; 
		block_ram[3291] = 24'b000000100000000010000000 ; 
		block_ram[3292] = 24'b000100000000011000000000 ; 
		block_ram[3293] = 24'b000000000010000100011000 ; 
		block_ram[3294] = 24'b000000011010000000100000 ; 
		block_ram[3295] = 24'b000000100000000010000100 ; 
		block_ram[3296] = 24'b100000000000001000000010 ; 
		block_ram[3297] = 24'b000000000010000100100100 ; 
		block_ram[3298] = 24'b100000000000001000000000 ; 
		block_ram[3299] = 24'b100000000000001000000001 ; 
		block_ram[3300] = 24'b000000000010000100100001 ; 
		block_ram[3301] = 24'b000000000010000100100000 ; 
		block_ram[3302] = 24'b100000000000001000000100 ; 
		block_ram[3303] = 24'b000000000010000100100010 ; 
		block_ram[3304] = 24'b000000001001010000000001 ; 
		block_ram[3305] = 24'b000000001001010000000000 ; 
		block_ram[3306] = 24'b100000000000001000001000 ; 
		block_ram[3307] = 24'b000000001001010000000010 ; 
		block_ram[3308] = 24'b000001100000100000000000 ; 
		block_ram[3309] = 24'b000000000010000100101000 ; 
		block_ram[3310] = 24'b000000011010000000010000 ; 
		block_ram[3311] = 24'b001100000100000000000000 ; 
		block_ram[3312] = 24'b000000000101000010000100 ; 
		block_ram[3313] = 24'b000100010000100000000000 ; 
		block_ram[3314] = 24'b100000000000001000010000 ; 
		block_ram[3315] = 24'b000000100000000010101000 ; 
		block_ram[3316] = 24'b000000000101000010000000 ; 
		block_ram[3317] = 24'b000000000010000100110000 ; 
		block_ram[3318] = 24'b000000000101000010000010 ; 
		block_ram[3319] = 24'b000001000000010001000000 ; 
		block_ram[3320] = 24'b001000000000000101000000 ; 
		block_ram[3321] = 24'b000000001001010000010000 ; 
		block_ram[3322] = 24'b000000011010000000000100 ; 
		block_ram[3323] = 24'b000000100000000010100000 ; 
		block_ram[3324] = 24'b000000000101000010001000 ; 
		block_ram[3325] = 24'b110010000000000000000000 ; 
		block_ram[3326] = 24'b000000011010000000000000 ; 
		block_ram[3327] = 24'b000000000001101100000000 ; 
		block_ram[3328] = 24'b000000000000110100000000 ; 
		block_ram[3329] = 24'b000000000000110100000001 ; 
		block_ram[3330] = 24'b000000000000110100000010 ; 
		block_ram[3331] = 24'b000100000001000000100000 ; 
		block_ram[3332] = 24'b000000000000110100000100 ; 
		block_ram[3333] = 24'b000000000010000011000000 ; 
		block_ram[3334] = 24'b000000001000001000010000 ; 
		block_ram[3335] = 24'b000000000010000011000010 ; 
		block_ram[3336] = 24'b000000000000110100001000 ; 
		block_ram[3337] = 24'b010010001000000000000000 ; 
		block_ram[3338] = 24'b100000010010000000000000 ; 
		block_ram[3339] = 24'b000000000100011010000000 ; 
		block_ram[3340] = 24'b000100100100000000000000 ; 
		block_ram[3341] = 24'b000000000010000011001000 ; 
		block_ram[3342] = 24'b000000001000001000011000 ; 
		block_ram[3343] = 24'b001001000000100000000000 ; 
		block_ram[3344] = 24'b000000000000110100010000 ; 
		block_ram[3345] = 24'b000001010100000000000000 ; 
		block_ram[3346] = 24'b000000001000001000000100 ; 
		block_ram[3347] = 24'b000000001000001000000101 ; 
		block_ram[3348] = 24'b000000001000001000000010 ; 
		block_ram[3349] = 24'b000000000010000011010000 ; 
		block_ram[3350] = 24'b000000001000001000000000 ; 
		block_ram[3351] = 24'b000000001000001000000001 ; 
		block_ram[3352] = 24'b001000000000000010100000 ; 
		block_ram[3353] = 24'b000000100000000101000010 ; 
		block_ram[3354] = 24'b000000001000001000001100 ; 
		block_ram[3355] = 24'b000000100000000101000000 ; 
		block_ram[3356] = 24'b000000001000001000001010 ; 
		block_ram[3357] = 24'b100000000001010000000000 ; 
		block_ram[3358] = 24'b000000001000001000001000 ; 
		block_ram[3359] = 24'b000000001000001000001001 ; 
		block_ram[3360] = 24'b000000000000110100100000 ; 
		block_ram[3361] = 24'b000100000001000000000010 ; 
		block_ram[3362] = 24'b000100000001000000000001 ; 
		block_ram[3363] = 24'b000100000001000000000000 ; 
		block_ram[3364] = 24'b110001000000000000000000 ; 
		block_ram[3365] = 24'b000000000010000011100000 ; 
		block_ram[3366] = 24'b000000001000001000110000 ; 
		block_ram[3367] = 24'b000100000001000000000100 ; 
		block_ram[3368] = 24'b001000000000000010010000 ; 
		block_ram[3369] = 24'b000000010000001100000100 ; 
		block_ram[3370] = 24'b000001001100000100000000 ; 
		block_ram[3371] = 24'b000100000001000000001000 ; 
		block_ram[3372] = 24'b000000001011100000000000 ; 
		block_ram[3373] = 24'b000000010000001100000000 ; 
		block_ram[3374] = 24'b000010000000010001000000 ; 
		block_ram[3375] = 24'b000000010000001100000010 ; 
		block_ram[3376] = 24'b001000000000000010001000 ; 
		block_ram[3377] = 24'b000001010100000000100000 ; 
		block_ram[3378] = 24'b000000001000001000100100 ; 
		block_ram[3379] = 24'b000100000001000000010000 ; 
		block_ram[3380] = 24'b000000000101000101000000 ; 
		block_ram[3381] = 24'b000010100000100000000000 ; 
		block_ram[3382] = 24'b000000001000001000100000 ; 
		block_ram[3383] = 24'b000000001000001000100001 ; 
		block_ram[3384] = 24'b001000000000000010000000 ; 
		block_ram[3385] = 24'b001000000000000010000001 ; 
		block_ram[3386] = 24'b001000000000000010000010 ; 
		block_ram[3387] = 24'b000000011000110000000000 ; 
		block_ram[3388] = 24'b001000000000000010000100 ; 
		block_ram[3389] = 24'b000000010000001100010000 ; 
		block_ram[3390] = 24'b000000001000001000101000 ; 
		block_ram[3391] = 24'b010000000110000000000000 ; 
		block_ram[3392] = 24'b000000000000110101000000 ; 
		block_ram[3393] = 24'b000000000010000010000100 ; 
		block_ram[3394] = 24'b011000000100000000000000 ; 
		block_ram[3395] = 24'b000000000010000010000110 ; 
		block_ram[3396] = 24'b000000000010000010000001 ; 
		block_ram[3397] = 24'b000000000010000010000000 ; 
		block_ram[3398] = 24'b000000000010000010000011 ; 
		block_ram[3399] = 24'b000000000010000010000010 ; 
		block_ram[3400] = 24'b000001000001001000000000 ; 
		block_ram[3401] = 24'b000000000010000010001100 ; 
		block_ram[3402] = 24'b000000100000000100010001 ; 
		block_ram[3403] = 24'b000000100000000100010000 ; 
		block_ram[3404] = 24'b000000000010000010001001 ; 
		block_ram[3405] = 24'b000000000010000010001000 ; 
		block_ram[3406] = 24'b000010000000010000100000 ; 
		block_ram[3407] = 24'b000000000010000010001010 ; 
		block_ram[3408] = 24'b100110000000000000000000 ; 
		block_ram[3409] = 24'b000000000010000010010100 ; 
		block_ram[3410] = 24'b000000001000001001000100 ; 
		block_ram[3411] = 24'b000000100000000100001000 ; 
		block_ram[3412] = 24'b000000000010000010010001 ; 
		block_ram[3413] = 24'b000000000010000010010000 ; 
		block_ram[3414] = 24'b000000001000001001000000 ; 
		block_ram[3415] = 24'b000000000010000010010010 ; 
		block_ram[3416] = 24'b000000001110010000000000 ; 
		block_ram[3417] = 24'b000000100000000100000010 ; 
		block_ram[3418] = 24'b000000100000000100000001 ; 
		block_ram[3419] = 24'b000000100000000100000000 ; 
		block_ram[3420] = 24'b010000010000100000000000 ; 
		block_ram[3421] = 24'b000000000010000010011000 ; 
		block_ram[3422] = 24'b000000001000001001001000 ; 
		block_ram[3423] = 24'b000000100000000100000100 ; 
		block_ram[3424] = 24'b000000111000000000000000 ; 
		block_ram[3425] = 24'b000000000010000010100100 ; 
		block_ram[3426] = 24'b000000111000000000000010 ; 
		block_ram[3427] = 24'b000100000001000001000000 ; 
		block_ram[3428] = 24'b000000000010000010100001 ; 
		block_ram[3429] = 24'b000000000010000010100000 ; 
		block_ram[3430] = 24'b000010000000010000001000 ; 
		block_ram[3431] = 24'b000000000010000010100010 ; 
		block_ram[3432] = 24'b000000111000000000001000 ; 
		block_ram[3433] = 24'b100000000100100000000000 ; 
		block_ram[3434] = 24'b000010000000010000000100 ; 
		block_ram[3435] = 24'b000000100000000100110000 ; 
		block_ram[3436] = 24'b000010000000010000000010 ; 
		block_ram[3437] = 24'b000000000010000010101000 ; 
		block_ram[3438] = 24'b000010000000010000000000 ; 
		block_ram[3439] = 24'b000010000000010000000001 ; 
		block_ram[3440] = 24'b000000000101000100000100 ; 
		block_ram[3441] = 24'b010000000000011000000000 ; 
		block_ram[3442] = 24'b000001000010100000000000 ; 
		block_ram[3443] = 24'b000000100000000100101000 ; 
		block_ram[3444] = 24'b000000000101000100000000 ; 
		block_ram[3445] = 24'b000000000010000010110000 ; 
		block_ram[3446] = 24'b000000000101000100000010 ; 
		block_ram[3447] = 24'b101000010000000000000000 ; 
		block_ram[3448] = 24'b001000000000000011000000 ; 
		block_ram[3449] = 24'b000000100000000100100010 ; 
		block_ram[3450] = 24'b000000100000000100100001 ; 
		block_ram[3451] = 24'b000000100000000100100000 ; 
		block_ram[3452] = 24'b000000000101000100001000 ; 
		block_ram[3453] = 24'b000101001000000000000000 ; 
		block_ram[3454] = 24'b000010000000010000010000 ; 
		block_ram[3455] = 24'b000000000001101010000000 ; 
		block_ram[3456] = 24'b000000000000110110000000 ; 
		block_ram[3457] = 24'b000000000010000001000100 ; 
		block_ram[3458] = 24'b000011100000000000000000 ; 
		block_ram[3459] = 24'b000000000010000001000110 ; 
		block_ram[3460] = 24'b000000000010000001000001 ; 
		block_ram[3461] = 24'b000000000010000001000000 ; 
		block_ram[3462] = 24'b000000000010000001000011 ; 
		block_ram[3463] = 24'b000000000010000001000010 ; 
		block_ram[3464] = 24'b001000000000000000110000 ; 
		block_ram[3465] = 24'b000000000010000001001100 ; 
		block_ram[3466] = 24'b000000000100011000000001 ; 
		block_ram[3467] = 24'b000000000100011000000000 ; 
		block_ram[3468] = 24'b000000000010000001001001 ; 
		block_ram[3469] = 24'b000000000010000001001000 ; 
		block_ram[3470] = 24'b010000000001000100000000 ; 
		block_ram[3471] = 24'b000000000010000001001010 ; 
		block_ram[3472] = 24'b001000000000000000101000 ; 
		block_ram[3473] = 24'b000000000010000001010100 ; 
		block_ram[3474] = 24'b000000001000001010000100 ; 
		block_ram[3475] = 24'b110000000000100000000000 ; 
		block_ram[3476] = 24'b000000000010000001010001 ; 
		block_ram[3477] = 24'b000000000010000001010000 ; 
		block_ram[3478] = 24'b000000001000001010000000 ; 
		block_ram[3479] = 24'b000000000010000001010010 ; 
		block_ram[3480] = 24'b001000000000000000100000 ; 
		block_ram[3481] = 24'b001000000000000000100001 ; 
		block_ram[3482] = 24'b001000000000000000100010 ; 
		block_ram[3483] = 24'b000000000100011000010000 ; 
		block_ram[3484] = 24'b001000000000000000100100 ; 
		block_ram[3485] = 24'b000000000010000001011000 ; 
		block_ram[3486] = 24'b000000001000001010001000 ; 
		block_ram[3487] = 24'b000110010000000000000000 ; 
		block_ram[3488] = 24'b001000000000000000011000 ; 
		block_ram[3489] = 24'b000000000010000001100100 ; 
		block_ram[3490] = 24'b000000010100100000000100 ; 
		block_ram[3491] = 24'b000100000001000010000000 ; 
		block_ram[3492] = 24'b000000000010000001100001 ; 
		block_ram[3493] = 24'b000000000010000001100000 ; 
		block_ram[3494] = 24'b000000010100100000000000 ; 
		block_ram[3495] = 24'b000000000010000001100010 ; 
		block_ram[3496] = 24'b001000000000000000010000 ; 
		block_ram[3497] = 24'b001000000000000000010001 ; 
		block_ram[3498] = 24'b001000000000000000010010 ; 
		block_ram[3499] = 24'b000000000100011000100000 ; 
		block_ram[3500] = 24'b001000000000000000010100 ; 
		block_ram[3501] = 24'b000000000010000001101000 ; 
		block_ram[3502] = 24'b000000010100100000001000 ; 
		block_ram[3503] = 24'b100000101000000000000000 ; 
		block_ram[3504] = 24'b001000000000000000001000 ; 
		block_ram[3505] = 24'b001000000000000000001001 ; 
		block_ram[3506] = 24'b001000000000000000001010 ; 
		block_ram[3507] = 24'b000000110010001000000000 ; 
		block_ram[3508] = 24'b001000000000000000001100 ; 
		block_ram[3509] = 24'b000000000010000001110000 ; 
		block_ram[3510] = 24'b000000001000001010100000 ; 
		block_ram[3511] = 24'b000001000000010100000000 ; 
		block_ram[3512] = 24'b001000000000000000000000 ; 
		block_ram[3513] = 24'b001000000000000000000001 ; 
		block_ram[3514] = 24'b001000000000000000000010 ; 
		block_ram[3515] = 24'b001000000000000000000011 ; 
		block_ram[3516] = 24'b001000000000000000000100 ; 
		block_ram[3517] = 24'b001000000000000000000101 ; 
		block_ram[3518] = 24'b001000000000000000000110 ; 
		block_ram[3519] = 24'b000000000001101001000000 ; 
		block_ram[3520] = 24'b000000000010000000000101 ; 
		block_ram[3521] = 24'b000000000010000000000100 ; 
		block_ram[3522] = 24'b000000000010000000000111 ; 
		block_ram[3523] = 24'b000000000010000000000110 ; 
		block_ram[3524] = 24'b000000000010000000000001 ; 
		block_ram[3525] = 24'b000000000010000000000000 ; 
		block_ram[3526] = 24'b000000000010000000000011 ; 
		block_ram[3527] = 24'b000000000010000000000010 ; 
		block_ram[3528] = 24'b000000000010000000001101 ; 
		block_ram[3529] = 24'b000000000010000000001100 ; 
		block_ram[3530] = 24'b000100001000100000000000 ; 
		block_ram[3531] = 24'b000000000010000000001110 ; 
		block_ram[3532] = 24'b000000000010000000001001 ; 
		block_ram[3533] = 24'b000000000010000000001000 ; 
		block_ram[3534] = 24'b000000000010000000001011 ; 
		block_ram[3535] = 24'b000000000010000000001010 ; 
		block_ram[3536] = 24'b000000000010000000010101 ; 
		block_ram[3537] = 24'b000000000010000000010100 ; 
		block_ram[3538] = 24'b000000010001010000000000 ; 
		block_ram[3539] = 24'b000000000010000000010110 ; 
		block_ram[3540] = 24'b000000000010000000010001 ; 
		block_ram[3541] = 24'b000000000010000000010000 ; 
		block_ram[3542] = 24'b000000000010000000010011 ; 
		block_ram[3543] = 24'b000000000010000000010010 ; 
		block_ram[3544] = 24'b001000000000000001100000 ; 
		block_ram[3545] = 24'b000000000010000000011100 ; 
		block_ram[3546] = 24'b000000010001010000001000 ; 
		block_ram[3547] = 24'b000000100000000110000000 ; 
		block_ram[3548] = 24'b000000000010000000011001 ; 
		block_ram[3549] = 24'b000000000010000000011000 ; 
		block_ram[3550] = 24'b100001000100000000000000 ; 
		block_ram[3551] = 24'b000000000001101000100000 ; 
		block_ram[3552] = 24'b000000000010000000100101 ; 
		block_ram[3553] = 24'b000000000010000000100100 ; 
		block_ram[3554] = 24'b100000000000001100000000 ; 
		block_ram[3555] = 24'b000000000010000000100110 ; 
		block_ram[3556] = 24'b000000000010000000100001 ; 
		block_ram[3557] = 24'b000000000010000000100000 ; 
		block_ram[3558] = 24'b000000000010000000100011 ; 
		block_ram[3559] = 24'b000000000010000000100010 ; 
		block_ram[3560] = 24'b001000000000000001010000 ; 
		block_ram[3561] = 24'b000000000010000000101100 ; 
		block_ram[3562] = 24'b000000100111000000000000 ; 
		block_ram[3563] = 24'b010001010000000000000000 ; 
		block_ram[3564] = 24'b000000000010000000101001 ; 
		block_ram[3565] = 24'b000000000010000000101000 ; 
		block_ram[3566] = 24'b000010000000010010000000 ; 
		block_ram[3567] = 24'b000000000001101000010000 ; 
		block_ram[3568] = 24'b001000000000000001001000 ; 
		block_ram[3569] = 24'b000000000010000000110100 ; 
		block_ram[3570] = 24'b000000010001010000100000 ; 
		block_ram[3571] = 24'b000010001100000000000000 ; 
		block_ram[3572] = 24'b000000000010000000110001 ; 
		block_ram[3573] = 24'b000000000010000000110000 ; 
		block_ram[3574] = 24'b010100100000000000000000 ; 
		block_ram[3575] = 24'b000000000001101000001000 ; 
		block_ram[3576] = 24'b001000000000000001000000 ; 
		block_ram[3577] = 24'b001000000000000001000001 ; 
		block_ram[3578] = 24'b001000000000000001000010 ; 
		block_ram[3579] = 24'b000000000001101000000100 ; 
		block_ram[3580] = 24'b001000000000000001000100 ; 
		block_ram[3581] = 24'b000000000001101000000010 ; 
		block_ram[3582] = 24'b000000000001101000000001 ; 
		block_ram[3583] = 24'b000000000001101000000000 ; 
		block_ram[3584] = 24'b000000000000111000000000 ; 
		block_ram[3585] = 24'b000000000000111000000001 ; 
		block_ram[3586] = 24'b000000000000111000000010 ; 
		block_ram[3587] = 24'b010001000010000000000000 ; 
		block_ram[3588] = 24'b000000000000111000000100 ; 
		block_ram[3589] = 24'b000000010000000000101000 ; 
		block_ram[3590] = 24'b000000001000000100010000 ; 
		block_ram[3591] = 24'b000000001000000100010001 ; 
		block_ram[3592] = 24'b000000000000111000001000 ; 
		block_ram[3593] = 24'b000000010000000000100100 ; 
		block_ram[3594] = 24'b001110000000000000000000 ; 
		block_ram[3595] = 24'b000000000100010110000000 ; 
		block_ram[3596] = 24'b000000010000000000100001 ; 
		block_ram[3597] = 24'b000000010000000000100000 ; 
		block_ram[3598] = 24'b000000000110100001000000 ; 
		block_ram[3599] = 24'b000000010000000000100010 ; 
		block_ram[3600] = 24'b000000000000111000010000 ; 
		block_ram[3601] = 24'b000010000001000010000000 ; 
		block_ram[3602] = 24'b000000001000000100000100 ; 
		block_ram[3603] = 24'b000000001000000100000101 ; 
		block_ram[3604] = 24'b000000001000000100000010 ; 
		block_ram[3605] = 24'b000000001000000100000011 ; 
		block_ram[3606] = 24'b000000001000000100000000 ; 
		block_ram[3607] = 24'b000000001000000100000001 ; 
		block_ram[3608] = 24'b110000000100000000000000 ; 
		block_ram[3609] = 24'b000000010000000000110100 ; 
		block_ram[3610] = 24'b000000000011010000100000 ; 
		block_ram[3611] = 24'b000000100000001001000000 ; 
		block_ram[3612] = 24'b000000001000000100001010 ; 
		block_ram[3613] = 24'b000000010000000000110000 ; 
		block_ram[3614] = 24'b000000001000000100001000 ; 
		block_ram[3615] = 24'b000000001000000100001001 ; 
		block_ram[3616] = 24'b000000000000111000100000 ; 
		block_ram[3617] = 24'b000000010000000000001100 ; 
		block_ram[3618] = 24'b100000000000000011000000 ; 
		block_ram[3619] = 24'b000000010000000000001110 ; 
		block_ram[3620] = 24'b000000010000000000001001 ; 
		block_ram[3621] = 24'b000000010000000000001000 ; 
		block_ram[3622] = 24'b000000001000000100110000 ; 
		block_ram[3623] = 24'b000000010000000000001010 ; 
		block_ram[3624] = 24'b000000010000000000000101 ; 
		block_ram[3625] = 24'b000000010000000000000100 ; 
		block_ram[3626] = 24'b000000000011010000010000 ; 
		block_ram[3627] = 24'b000000010000000000000110 ; 
		block_ram[3628] = 24'b000000010000000000000001 ; 
		block_ram[3629] = 24'b000000010000000000000000 ; 
		block_ram[3630] = 24'b000000010000000000000011 ; 
		block_ram[3631] = 24'b000000010000000000000010 ; 
		block_ram[3632] = 24'b000101100000000000000000 ; 
		block_ram[3633] = 24'b000000010000000000011100 ; 
		block_ram[3634] = 24'b000000000011010000001000 ; 
		block_ram[3635] = 24'b001000000100100000000000 ; 
		block_ram[3636] = 24'b000000000101001001000000 ; 
		block_ram[3637] = 24'b000000010000000000011000 ; 
		block_ram[3638] = 24'b000000001000000100100000 ; 
		block_ram[3639] = 24'b000000001000000100100001 ; 
		block_ram[3640] = 24'b000000000011010000000010 ; 
		block_ram[3641] = 24'b000000010000000000010100 ; 
		block_ram[3642] = 24'b000000000011010000000000 ; 
		block_ram[3643] = 24'b000000000011010000000001 ; 
		block_ram[3644] = 24'b000000010000000000010001 ; 
		block_ram[3645] = 24'b000000010000000000010000 ; 
		block_ram[3646] = 24'b000000000011010000000100 ; 
		block_ram[3647] = 24'b000000010000000000010010 ; 
		block_ram[3648] = 24'b000000000000111001000000 ; 
		block_ram[3649] = 24'b000100001100000000000000 ; 
		block_ram[3650] = 24'b100000000000000010100000 ; 
		block_ram[3651] = 24'b000000100000001000011000 ; 
		block_ram[3652] = 24'b010010100000000000000000 ; 
		block_ram[3653] = 24'b000000000010001110000000 ; 
		block_ram[3654] = 24'b000000000110100000001000 ; 
		block_ram[3655] = 24'b001000000001010000000000 ; 
		block_ram[3656] = 24'b000001000001000100000000 ; 
		block_ram[3657] = 24'b000000010000000001100100 ; 
		block_ram[3658] = 24'b000000000110100000000100 ; 
		block_ram[3659] = 24'b000000100000001000010000 ; 
		block_ram[3660] = 24'b000000000110100000000010 ; 
		block_ram[3661] = 24'b000000010000000001100000 ; 
		block_ram[3662] = 24'b000000000110100000000000 ; 
		block_ram[3663] = 24'b000000000110100000000001 ; 
		block_ram[3664] = 24'b001000010010000000000000 ; 
		block_ram[3665] = 24'b000000100000001000001010 ; 
		block_ram[3666] = 24'b000000001000000101000100 ; 
		block_ram[3667] = 24'b000000100000001000001000 ; 
		block_ram[3668] = 24'b000000000101001000100000 ; 
		block_ram[3669] = 24'b100001000000100000000000 ; 
		block_ram[3670] = 24'b000000001000000101000000 ; 
		block_ram[3671] = 24'b000000001000000101000001 ; 
		block_ram[3672] = 24'b000000100000001000000011 ; 
		block_ram[3673] = 24'b000000100000001000000010 ; 
		block_ram[3674] = 24'b000000100000001000000001 ; 
		block_ram[3675] = 24'b000000100000001000000000 ; 
		block_ram[3676] = 24'b000100000000010010000000 ; 
		block_ram[3677] = 24'b000000010000000001110000 ; 
		block_ram[3678] = 24'b000000000110100000010000 ; 
		block_ram[3679] = 24'b000000100000001000000100 ; 
		block_ram[3680] = 24'b100000000000000010000010 ; 
		block_ram[3681] = 24'b000000010000000001001100 ; 
		block_ram[3682] = 24'b100000000000000010000000 ; 
		block_ram[3683] = 24'b100000000000000010000001 ; 
		block_ram[3684] = 24'b000000000101001000010000 ; 
		block_ram[3685] = 24'b000000010000000001001000 ; 
		block_ram[3686] = 24'b100000000000000010000100 ; 
		block_ram[3687] = 24'b000000010000000001001010 ; 
		block_ram[3688] = 24'b000000010000000001000101 ; 
		block_ram[3689] = 24'b000000010000000001000100 ; 
		block_ram[3690] = 24'b100000000000000010001000 ; 
		block_ram[3691] = 24'b000000010000000001000110 ; 
		block_ram[3692] = 24'b000000010000000001000001 ; 
		block_ram[3693] = 24'b000000010000000001000000 ; 
		block_ram[3694] = 24'b000000000110100000100000 ; 
		block_ram[3695] = 24'b000000010000000001000010 ; 
		block_ram[3696] = 24'b000000000101001000000100 ; 
		block_ram[3697] = 24'b010000000000010100000000 ; 
		block_ram[3698] = 24'b100000000000000010010000 ; 
		block_ram[3699] = 24'b000000100000001000101000 ; 
		block_ram[3700] = 24'b000000000101001000000000 ; 
		block_ram[3701] = 24'b000000000101001000000001 ; 
		block_ram[3702] = 24'b000000000101001000000010 ; 
		block_ram[3703] = 24'b000110000010000000000000 ; 
		block_ram[3704] = 24'b000010001000100000000000 ; 
		block_ram[3705] = 24'b000000010000000001010100 ; 
		block_ram[3706] = 24'b000000000011010001000000 ; 
		block_ram[3707] = 24'b000000100000001000100000 ; 
		block_ram[3708] = 24'b000000000101001000001000 ; 
		block_ram[3709] = 24'b000000010000000001010000 ; 
		block_ram[3710] = 24'b011001000000000000000000 ; 
		block_ram[3711] = 24'b000000000001100110000000 ; 
		block_ram[3712] = 24'b000000000000111010000000 ; 
		block_ram[3713] = 24'b000010000001000000010000 ; 
		block_ram[3714] = 24'b100000000000000001100000 ; 
		block_ram[3715] = 24'b000000000100010100001000 ; 
		block_ram[3716] = 24'b001001000100000000000000 ; 
		block_ram[3717] = 24'b000000000010001101000000 ; 
		block_ram[3718] = 24'b000000001000000110010000 ; 
		block_ram[3719] = 24'b000100100000100000000000 ; 
		block_ram[3720] = 24'b000000101010000000000000 ; 
		block_ram[3721] = 24'b000000000100010100000010 ; 
		block_ram[3722] = 24'b000000000100010100000001 ; 
		block_ram[3723] = 24'b000000000100010100000000 ; 
		block_ram[3724] = 24'b000000010000000010100001 ; 
		block_ram[3725] = 24'b000000010000000010100000 ; 
		block_ram[3726] = 24'b010000000001001000000000 ; 
		block_ram[3727] = 24'b000000000100010100000100 ; 
		block_ram[3728] = 24'b000010000001000000000001 ; 
		block_ram[3729] = 24'b000010000001000000000000 ; 
		block_ram[3730] = 24'b000000001000000110000100 ; 
		block_ram[3731] = 24'b000010000001000000000010 ; 
		block_ram[3732] = 24'b000000001000000110000010 ; 
		block_ram[3733] = 24'b000010000001000000000100 ; 
		block_ram[3734] = 24'b000000001000000110000000 ; 
		block_ram[3735] = 24'b000000001000000110000001 ; 
		block_ram[3736] = 24'b000000101010000000010000 ; 
		block_ram[3737] = 24'b000010000001000000001000 ; 
		block_ram[3738] = 24'b000001010000100000000000 ; 
		block_ram[3739] = 24'b000000000100010100010000 ; 
		block_ram[3740] = 24'b000100000000010001000000 ; 
		block_ram[3741] = 24'b000000001100101000000000 ; 
		block_ram[3742] = 24'b000000001000000110001000 ; 
		block_ram[3743] = 24'b101000000010000000000000 ; 
		block_ram[3744] = 24'b100000000000000001000010 ; 
		block_ram[3745] = 24'b000000010000000010001100 ; 
		block_ram[3746] = 24'b100000000000000001000000 ; 
		block_ram[3747] = 24'b100000000000000001000001 ; 
		block_ram[3748] = 24'b000000010000000010001001 ; 
		block_ram[3749] = 24'b000000010000000010001000 ; 
		block_ram[3750] = 24'b100000000000000001000100 ; 
		block_ram[3751] = 24'b000000001111000000000000 ; 
		block_ram[3752] = 24'b000000010000000010000101 ; 
		block_ram[3753] = 24'b000000010000000010000100 ; 
		block_ram[3754] = 24'b100000000000000001001000 ; 
		block_ram[3755] = 24'b000000000100010100100000 ; 
		block_ram[3756] = 24'b000000010000000010000001 ; 
		block_ram[3757] = 24'b000000010000000010000000 ; 
		block_ram[3758] = 24'b000000010000000010000011 ; 
		block_ram[3759] = 24'b000000010000000010000010 ; 
		block_ram[3760] = 24'b000000011100010000000000 ; 
		block_ram[3761] = 24'b000010000001000000100000 ; 
		block_ram[3762] = 24'b100000000000000001010000 ; 
		block_ram[3763] = 24'b000000110010000100000000 ; 
		block_ram[3764] = 24'b010000000010100000000000 ; 
		block_ram[3765] = 24'b000000010000000010011000 ; 
		block_ram[3766] = 24'b000000001000000110100000 ; 
		block_ram[3767] = 24'b000001000000011000000000 ; 
		block_ram[3768] = 24'b001000000000001100000000 ; 
		block_ram[3769] = 24'b000000010000000010010100 ; 
		block_ram[3770] = 24'b000000000011010010000000 ; 
		block_ram[3771] = 24'b010100001000000000000000 ; 
		block_ram[3772] = 24'b000000010000000010010001 ; 
		block_ram[3773] = 24'b000000010000000010010000 ; 
		block_ram[3774] = 24'b000010100100000000000000 ; 
		block_ram[3775] = 24'b000000000001100101000000 ; 
		block_ram[3776] = 24'b100000000000000000100010 ; 
		block_ram[3777] = 24'b000000000010001100000100 ; 
		block_ram[3778] = 24'b100000000000000000100000 ; 
		block_ram[3779] = 24'b100000000000000000100001 ; 
		block_ram[3780] = 24'b000000000010001100000001 ; 
		block_ram[3781] = 24'b000000000010001100000000 ; 
		block_ram[3782] = 24'b100000000000000000100100 ; 
		block_ram[3783] = 24'b000000000010001100000010 ; 
		block_ram[3784] = 24'b000000101010000001000000 ; 
		block_ram[3785] = 24'b011000000000100000000000 ; 
		block_ram[3786] = 24'b100000000000000000101000 ; 
		block_ram[3787] = 24'b000000000100010101000000 ; 
		block_ram[3788] = 24'b000100000000010000010000 ; 
		block_ram[3789] = 24'b000000000010001100001000 ; 
		block_ram[3790] = 24'b000000000110100010000000 ; 
		block_ram[3791] = 24'b000011001000000000000000 ; 
		block_ram[3792] = 24'b000000100100100100000000 ; 
		block_ram[3793] = 24'b000010000001000001000000 ; 
		block_ram[3794] = 24'b100000000000000000110000 ; 
		block_ram[3795] = 24'b000000001010110000000000 ; 
		block_ram[3796] = 24'b000100000000010000001000 ; 
		block_ram[3797] = 24'b000000000010001100010000 ; 
		block_ram[3798] = 24'b000000001000000111000000 ; 
		block_ram[3799] = 24'b010000010100000000000000 ; 
		block_ram[3800] = 24'b000100000000010000000100 ; 
		block_ram[3801] = 24'b000000100000001010000010 ; 
		block_ram[3802] = 24'b000000100000001010000001 ; 
		block_ram[3803] = 24'b000000100000001010000000 ; 
		block_ram[3804] = 24'b000100000000010000000000 ; 
		block_ram[3805] = 24'b000100000000010000000001 ; 
		block_ram[3806] = 24'b000100000000010000000010 ; 
		block_ram[3807] = 24'b000000000001100100100000 ; 
		block_ram[3808] = 24'b100000000000000000000010 ; 
		block_ram[3809] = 24'b100000000000000000000011 ; 
		block_ram[3810] = 24'b100000000000000000000000 ; 
		block_ram[3811] = 24'b100000000000000000000001 ; 
		block_ram[3812] = 24'b100000000000000000000110 ; 
		block_ram[3813] = 24'b000000000010001100100000 ; 
		block_ram[3814] = 24'b100000000000000000000100 ; 
		block_ram[3815] = 24'b100000000000000000000101 ; 
		block_ram[3816] = 24'b100000000000000000001010 ; 
		block_ram[3817] = 24'b000000001001011000000000 ; 
		block_ram[3818] = 24'b100000000000000000001000 ; 
		block_ram[3819] = 24'b100000000000000000001001 ; 
		block_ram[3820] = 24'b000000010000000011000001 ; 
		block_ram[3821] = 24'b000000010000000011000000 ; 
		block_ram[3822] = 24'b100000000000000000001100 ; 
		block_ram[3823] = 24'b000000000001100100010000 ; 
		block_ram[3824] = 24'b100000000000000000010010 ; 
		block_ram[3825] = 24'b000001000110000000001000 ; 
		block_ram[3826] = 24'b100000000000000000010000 ; 
		block_ram[3827] = 24'b100000000000000000010001 ; 
		block_ram[3828] = 24'b000000000101001010000000 ; 
		block_ram[3829] = 24'b001000101000000000000000 ; 
		block_ram[3830] = 24'b100000000000000000010100 ; 
		block_ram[3831] = 24'b000000000001100100001000 ; 
		block_ram[3832] = 24'b000001000110000000000001 ; 
		block_ram[3833] = 24'b000001000110000000000000 ; 
		block_ram[3834] = 24'b100000000000000000011000 ; 
		block_ram[3835] = 24'b000000000001100100000100 ; 
		block_ram[3836] = 24'b000100000000010000100000 ; 
		block_ram[3837] = 24'b000000000001100100000010 ; 
		block_ram[3838] = 24'b000000000001100100000001 ; 
		block_ram[3839] = 24'b000000000001100100000000 ; 
		block_ram[3840] = 24'b000000000000111100000000 ; 
		block_ram[3841] = 24'b101000100000000000000000 ; 
		block_ram[3842] = 24'b000000001000000000010100 ; 
		block_ram[3843] = 24'b000000000100010010001000 ; 
		block_ram[3844] = 24'b000000001000000000010010 ; 
		block_ram[3845] = 24'b000000000010001011000000 ; 
		block_ram[3846] = 24'b000000001000000000010000 ; 
		block_ram[3847] = 24'b000000001000000000010001 ; 
		block_ram[3848] = 24'b000001000001000001000000 ; 
		block_ram[3849] = 24'b000000000100010010000010 ; 
		block_ram[3850] = 24'b000000000100010010000001 ; 
		block_ram[3851] = 24'b000000000100010010000000 ; 
		block_ram[3852] = 24'b000000001000000000011010 ; 
		block_ram[3853] = 24'b000000010000000100100000 ; 
		block_ram[3854] = 24'b000000001000000000011000 ; 
		block_ram[3855] = 24'b000000000100010010000100 ; 
		block_ram[3856] = 24'b000000001000000000000110 ; 
		block_ram[3857] = 24'b000000001000000000000111 ; 
		block_ram[3858] = 24'b000000001000000000000100 ; 
		block_ram[3859] = 24'b000000001000000000000101 ; 
		block_ram[3860] = 24'b000000001000000000000010 ; 
		block_ram[3861] = 24'b000000001000000000000011 ; 
		block_ram[3862] = 24'b000000001000000000000000 ; 
		block_ram[3863] = 24'b000000001000000000000001 ; 
		block_ram[3864] = 24'b000000001000000000001110 ; 
		block_ram[3865] = 24'b000100000010100000000000 ; 
		block_ram[3866] = 24'b000000001000000000001100 ; 
		block_ram[3867] = 24'b000000000100010010010000 ; 
		block_ram[3868] = 24'b000000001000000000001010 ; 
		block_ram[3869] = 24'b000000001000000000001011 ; 
		block_ram[3870] = 24'b000000001000000000001000 ; 
		block_ram[3871] = 24'b000000001000000000001001 ; 
		block_ram[3872] = 24'b000010000110000000000000 ; 
		block_ram[3873] = 24'b000000010000000100001100 ; 
		block_ram[3874] = 24'b000000001000000000110100 ; 
		block_ram[3875] = 24'b000100000001001000000000 ; 
		block_ram[3876] = 24'b000000001000000000110010 ; 
		block_ram[3877] = 24'b000000010000000100001000 ; 
		block_ram[3878] = 24'b000000001000000000110000 ; 
		block_ram[3879] = 24'b000000001000000000110001 ; 
		block_ram[3880] = 24'b000000010000000100000101 ; 
		block_ram[3881] = 24'b000000010000000100000100 ; 
		block_ram[3882] = 24'b010000100000100000000000 ; 
		block_ram[3883] = 24'b000000000100010010100000 ; 
		block_ram[3884] = 24'b000000010000000100000001 ; 
		block_ram[3885] = 24'b000000010000000100000000 ; 
		block_ram[3886] = 24'b000000001000000000111000 ; 
		block_ram[3887] = 24'b000000010000000100000010 ; 
		block_ram[3888] = 24'b000000001000000000100110 ; 
		block_ram[3889] = 24'b010000000000010001000000 ; 
		block_ram[3890] = 24'b000000001000000000100100 ; 
		block_ram[3891] = 24'b000000001000000000100101 ; 
		block_ram[3892] = 24'b000000001000000000100010 ; 
		block_ram[3893] = 24'b000000001000000000100011 ; 
		block_ram[3894] = 24'b000000001000000000100000 ; 
		block_ram[3895] = 24'b000000001000000000100001 ; 
		block_ram[3896] = 24'b001000000000001010000000 ; 
		block_ram[3897] = 24'b000000010000000100010100 ; 
		block_ram[3898] = 24'b000000000011010100000000 ; 
		block_ram[3899] = 24'b100011000000000000000000 ; 
		block_ram[3900] = 24'b000000001000000000101010 ; 
		block_ram[3901] = 24'b000000010000000100010000 ; 
		block_ram[3902] = 24'b000000001000000000101000 ; 
		block_ram[3903] = 24'b000000000001100011000000 ; 
		block_ram[3904] = 24'b000001000001000000001000 ; 
		block_ram[3905] = 24'b000000000010001010000100 ; 
		block_ram[3906] = 24'b000000001000000001010100 ; 
		block_ram[3907] = 24'b000010010000100000000000 ; 
		block_ram[3908] = 24'b000000000010001010000001 ; 
		block_ram[3909] = 24'b000000000010001010000000 ; 
		block_ram[3910] = 24'b000000001000000001010000 ; 
		block_ram[3911] = 24'b000000000010001010000010 ; 
		block_ram[3912] = 24'b000001000001000000000000 ; 
		block_ram[3913] = 24'b000001000001000000000001 ; 
		block_ram[3914] = 24'b000001000001000000000010 ; 
		block_ram[3915] = 24'b000000000100010011000000 ; 
		block_ram[3916] = 24'b000001000001000000000100 ; 
		block_ram[3917] = 24'b000000000010001010001000 ; 
		block_ram[3918] = 24'b000000000110100100000000 ; 
		block_ram[3919] = 24'b110100000000000000000000 ; 
		block_ram[3920] = 24'b000000001000000001000110 ; 
		block_ram[3921] = 24'b010000000000010000100000 ; 
		block_ram[3922] = 24'b000000001000000001000100 ; 
		block_ram[3923] = 24'b000000001000000001000101 ; 
		block_ram[3924] = 24'b000000001000000001000010 ; 
		block_ram[3925] = 24'b000000000010001010010000 ; 
		block_ram[3926] = 24'b000000001000000001000000 ; 
		block_ram[3927] = 24'b000000001000000001000001 ; 
		block_ram[3928] = 24'b000001000001000000010000 ; 
		block_ram[3929] = 24'b000000100000001100000010 ; 
		block_ram[3930] = 24'b000000001000000001001100 ; 
		block_ram[3931] = 24'b000000100000001100000000 ; 
		block_ram[3932] = 24'b000000001000000001001010 ; 
		block_ram[3933] = 24'b001010000100000000000000 ; 
		block_ram[3934] = 24'b000000001000000001001000 ; 
		block_ram[3935] = 24'b000000000001100010100000 ; 
		block_ram[3936] = 24'b000000111000001000000000 ; 
		block_ram[3937] = 24'b010000000000010000010000 ; 
		block_ram[3938] = 24'b100000000000000110000000 ; 
		block_ram[3939] = 24'b000001100100000000000100 ; 
		block_ram[3940] = 24'b001100000000100000000000 ; 
		block_ram[3941] = 24'b000000000010001010100000 ; 
		block_ram[3942] = 24'b000000001000000001110000 ; 
		block_ram[3943] = 24'b000001100100000000000000 ; 
		block_ram[3944] = 24'b000001000001000000100000 ; 
		block_ram[3945] = 24'b000000010000000101000100 ; 
		block_ram[3946] = 24'b000001000001000000100010 ; 
		block_ram[3947] = 24'b001000001010000000000000 ; 
		block_ram[3948] = 24'b000000010000000101000001 ; 
		block_ram[3949] = 24'b000000010000000101000000 ; 
		block_ram[3950] = 24'b000010000000011000000000 ; 
		block_ram[3951] = 24'b000000000001100010010000 ; 
		block_ram[3952] = 24'b010000000000010000000001 ; 
		block_ram[3953] = 24'b010000000000010000000000 ; 
		block_ram[3954] = 24'b000000001000000001100100 ; 
		block_ram[3955] = 24'b010000000000010000000010 ; 
		block_ram[3956] = 24'b000000000101001100000000 ; 
		block_ram[3957] = 24'b010000000000010000000100 ; 
		block_ram[3958] = 24'b000000001000000001100000 ; 
		block_ram[3959] = 24'b000000000001100010001000 ; 
		block_ram[3960] = 24'b000001000001000000110000 ; 
		block_ram[3961] = 24'b010000000000010000001000 ; 
		block_ram[3962] = 24'b000100010100000000000000 ; 
		block_ram[3963] = 24'b000000000001100010000100 ; 
		block_ram[3964] = 24'b100000100010000000000000 ; 
		block_ram[3965] = 24'b000000000001100010000010 ; 
		block_ram[3966] = 24'b000000000001100010000001 ; 
		block_ram[3967] = 24'b000000000001100010000000 ; 
		block_ram[3968] = 24'b010100010000000000000000 ; 
		block_ram[3969] = 24'b000000000010001001000100 ; 
		block_ram[3970] = 24'b000000000100010000001001 ; 
		block_ram[3971] = 24'b000000000100010000001000 ; 
		block_ram[3972] = 24'b000000000010001001000001 ; 
		block_ram[3973] = 24'b000000000010001001000000 ; 
		block_ram[3974] = 24'b000000001000000010010000 ; 
		block_ram[3975] = 24'b000000000010001001000010 ; 
		block_ram[3976] = 24'b000000000100010000000011 ; 
		block_ram[3977] = 24'b000000000100010000000010 ; 
		block_ram[3978] = 24'b000000000100010000000001 ; 
		block_ram[3979] = 24'b000000000100010000000000 ; 
		block_ram[3980] = 24'b100010000000100000000000 ; 
		block_ram[3981] = 24'b000000000010001001001000 ; 
		block_ram[3982] = 24'b000000000100010000000101 ; 
		block_ram[3983] = 24'b000000000100010000000100 ; 
		block_ram[3984] = 24'b000000001000000010000110 ; 
		block_ram[3985] = 24'b000010000001000100000000 ; 
		block_ram[3986] = 24'b000000001000000010000100 ; 
		block_ram[3987] = 24'b000000000100010000011000 ; 
		block_ram[3988] = 24'b000000001000000010000010 ; 
		block_ram[3989] = 24'b000000000010001001010000 ; 
		block_ram[3990] = 24'b000000001000000010000000 ; 
		block_ram[3991] = 24'b000000001000000010000001 ; 
		block_ram[3992] = 24'b001000000000001000100000 ; 
		block_ram[3993] = 24'b000000000100010000010010 ; 
		block_ram[3994] = 24'b000000000100010000010001 ; 
		block_ram[3995] = 24'b000000000100010000010000 ; 
		block_ram[3996] = 24'b000000001000000010001010 ; 
		block_ram[3997] = 24'b010001100000000000000000 ; 
		block_ram[3998] = 24'b000000001000000010001000 ; 
		block_ram[3999] = 24'b000000000001100001100000 ; 
		block_ram[4000] = 24'b000000100001010000000100 ; 
		block_ram[4001] = 24'b000001001000100000000000 ; 
		block_ram[4002] = 24'b100000000000000101000000 ; 
		block_ram[4003] = 24'b000000000100010000101000 ; 
		block_ram[4004] = 24'b000000100001010000000000 ; 
		block_ram[4005] = 24'b000000000010001001100000 ; 
		block_ram[4006] = 24'b000000001000000010110000 ; 
		block_ram[4007] = 24'b011010000000000000000000 ; 
		block_ram[4008] = 24'b001000000000001000010000 ; 
		block_ram[4009] = 24'b000000000100010000100010 ; 
		block_ram[4010] = 24'b000000000100010000100001 ; 
		block_ram[4011] = 24'b000000000100010000100000 ; 
		block_ram[4012] = 24'b000000010000000110000001 ; 
		block_ram[4013] = 24'b000000010000000110000000 ; 
		block_ram[4014] = 24'b000101000010000000000000 ; 
		block_ram[4015] = 24'b000000000001100001010000 ; 
		block_ram[4016] = 24'b001000000000001000001000 ; 
		block_ram[4017] = 24'b000000110010000000000010 ; 
		block_ram[4018] = 24'b000000001000000010100100 ; 
		block_ram[4019] = 24'b000000110010000000000000 ; 
		block_ram[4020] = 24'b000000001000000010100010 ; 
		block_ram[4021] = 24'b100100000100000000000000 ; 
		block_ram[4022] = 24'b000000001000000010100000 ; 
		block_ram[4023] = 24'b000000000001100001001000 ; 
		block_ram[4024] = 24'b001000000000001000000000 ; 
		block_ram[4025] = 24'b001000000000001000000001 ; 
		block_ram[4026] = 24'b001000000000001000000010 ; 
		block_ram[4027] = 24'b000000000001100001000100 ; 
		block_ram[4028] = 24'b001000000000001000000100 ; 
		block_ram[4029] = 24'b000000000001100001000010 ; 
		block_ram[4030] = 24'b000000000001100001000001 ; 
		block_ram[4031] = 24'b000000000001100001000000 ; 
		block_ram[4032] = 24'b000000000010001000000101 ; 
		block_ram[4033] = 24'b000000000010001000000100 ; 
		block_ram[4034] = 24'b100000000000000100100000 ; 
		block_ram[4035] = 24'b000000000010001000000110 ; 
		block_ram[4036] = 24'b000000000010001000000001 ; 
		block_ram[4037] = 24'b000000000010001000000000 ; 
		block_ram[4038] = 24'b000000000010001000000011 ; 
		block_ram[4039] = 24'b000000000010001000000010 ; 
		block_ram[4040] = 24'b000001000001000010000000 ; 
		block_ram[4041] = 24'b000000000010001000001100 ; 
		block_ram[4042] = 24'b000000000100010001000001 ; 
		block_ram[4043] = 24'b000000000100010001000000 ; 
		block_ram[4044] = 24'b000000000010001000001001 ; 
		block_ram[4045] = 24'b000000000010001000001000 ; 
		block_ram[4046] = 24'b001000110000000000000000 ; 
		block_ram[4047] = 24'b000000000001100000110000 ; 
		block_ram[4048] = 24'b000000100100100000000000 ; 
		block_ram[4049] = 24'b000000000010001000010100 ; 
		block_ram[4050] = 24'b000000001000000011000100 ; 
		block_ram[4051] = 24'b001101000000000000000000 ; 
		block_ram[4052] = 24'b000000000010001000010001 ; 
		block_ram[4053] = 24'b000000000010001000010000 ; 
		block_ram[4054] = 24'b000000001000000011000000 ; 
		block_ram[4055] = 24'b000000000001100000101000 ; 
		block_ram[4056] = 24'b000000100100100000001000 ; 
		block_ram[4057] = 24'b100000011000000000000000 ; 
		block_ram[4058] = 24'b010010000010000000000000 ; 
		block_ram[4059] = 24'b000000000001100000100100 ; 
		block_ram[4060] = 24'b000100000000010100000000 ; 
		block_ram[4061] = 24'b000000000001100000100010 ; 
		block_ram[4062] = 24'b000000000001100000100001 ; 
		block_ram[4063] = 24'b000000000001100000100000 ; 
		block_ram[4064] = 24'b100000000000000100000010 ; 
		block_ram[4065] = 24'b000000000010001000100100 ; 
		block_ram[4066] = 24'b100000000000000100000000 ; 
		block_ram[4067] = 24'b100000000000000100000001 ; 
		block_ram[4068] = 24'b000000000010001000100001 ; 
		block_ram[4069] = 24'b000000000010001000100000 ; 
		block_ram[4070] = 24'b100000000000000100000100 ; 
		block_ram[4071] = 24'b000000000001100000011000 ; 
		block_ram[4072] = 24'b000000010010110000000000 ; 
		block_ram[4073] = 24'b000110100000000000000000 ; 
		block_ram[4074] = 24'b100000000000000100001000 ; 
		block_ram[4075] = 24'b000000000001100000010100 ; 
		block_ram[4076] = 24'b010000001100000000000000 ; 
		block_ram[4077] = 24'b000000000001100000010010 ; 
		block_ram[4078] = 24'b000000000001100000010001 ; 
		block_ram[4079] = 24'b000000000001100000010000 ; 
		block_ram[4080] = 24'b000000100100100000100000 ; 
		block_ram[4081] = 24'b010000000000010010000000 ; 
		block_ram[4082] = 24'b100000000000000100010000 ; 
		block_ram[4083] = 24'b000000000001100000001100 ; 
		block_ram[4084] = 24'b000011010000000000000000 ; 
		block_ram[4085] = 24'b000000000001100000001010 ; 
		block_ram[4086] = 24'b000000000001100000001001 ; 
		block_ram[4087] = 24'b000000000001100000001000 ; 
		block_ram[4088] = 24'b001000000000001001000000 ; 
		block_ram[4089] = 24'b000000000001100000000110 ; 
		block_ram[4090] = 24'b000000000001100000000101 ; 
		block_ram[4091] = 24'b000000000001100000000100 ; 
		block_ram[4092] = 24'b000000000001100000000011 ; 
		block_ram[4093] = 24'b000000000001100000000010 ; 
		block_ram[4094] = 24'b000000000001100000000001 ; 
		block_ram[4095] = 24'b000000000001100000000000 ; 
	end

   always @(posedge clk)
	begin
      output_reg <= block_ram[address];
	end



endmodule
